module pixel_itr(
    input wire clk,
    input wire pix_clk,
    input wire rst,
    output wire [9:0] pix_x,
    output wire [9:0] pix_y,
    output wire h_sync,
    output wire v_sync,
    output wire draw_active,
    output wire screen_end,
    output wire draw_end
    );
	 
	// FOR 800 X 600
    // parameter h_sync_strt = 56;          
    // parameter h_sync_end  = 56 + 120;         
    // parameter v_sync_strt = 600 + 37;        
    // parameter v_sync_end  = 600 + 37 + 6;   
    // parameter h_draw_min  = 56 + 120 + 64;   
    // parameter v_draw_max  = 600 - 1;            
    // parameter h_max = 1040;           
    // parameter v_max = 666 - 1;
	 
	// FOR 640 X 480
    parameter h_sync_strt = 16;          
    parameter h_sync_end  = 16 + 96;         
    parameter v_sync_strt = 480 + 10;        
    parameter v_sync_end  = 480 + 10 + 2;   
    parameter h_draw_min  = 16 + 96 + 48;   
    parameter v_draw_max  = 480 - 1;            
    parameter h_max = 800;           
    parameter v_max = 525 - 1;

    reg [9:0] h_pos=0;
	 reg [9:0] v_pos=0; 
	
    // --------------- SYNC SIGNALS BLOCK ---------------
    assign h_sync = (h_pos >= h_sync_strt && h_pos < h_sync_end) ? 0 : 1;
    assign v_sync = (v_pos >= v_sync_strt && v_pos < v_sync_end) ? 0 : 1;
    // --------------------------------------------------
		
	// -------------- PIXEL POSITION BLOCK --------------
    // assign pix_x = (h_pos >= h_draw_min) ? h_pos : 0;        
    assign pix_x = (h_pos >= h_draw_min) ? h_pos - h_draw_min : 0;        
	 assign pix_y = (v_pos <= v_draw_max) ? v_pos : v_draw_max;        
    // --------------------------------------------------

    // -------- BLANKING / DRAWING PERIOD BLOCK ---------
    assign draw_active = (h_pos < h_draw_min | v_pos > v_draw_max) ? 0 : 1;
    // --------------------------------------------------

    // ----------------- LIMITS BLOCK -------------------
    assign screen_end = (h_pos == h_max & v_pos == v_max);
    assign draw_end = (h_pos == h_max & v_pos == v_draw_max);
    // --------------------------------------------------
    
    // ------------------ MAIN BLOCK --------------------
    always @ (posedge clk) begin
        if (rst) begin
            h_pos <= 0; 
            v_pos <= 0;
        end

        if(pix_clk) begin
            if (h_pos < h_max) begin
                h_pos <= h_pos + 1; 
            end
            else begin
                h_pos <= 0;
                v_pos <= v_pos + 1;
            end

            if (v_pos == v_max) begin
                    v_pos <= 0;
            end
        end
    end
    // --------------------------------------------------

endmodule

//////////////////////////////////////////////////////////////////////////////////

module screen_design(
	input clk,
	input rst,
	output h_sync,
	output v_sync,
	output r_out,
	output g_out,
	output b_out
);

//---------------GENERATING PIXEL CLOCK----------------------
reg count = 0, pix_clk = 0;

always @(posedge clk) begin
	
	if (rst == 1) begin
		count <= 0;
		pix_clk <= 0;
	end 
	if (count == 1) begin
		pix_clk <= 1;
		count <= 0;
	end 
	else begin
		pix_clk <= 0;
		count <= count + 1;

	end
end

//-----------------------------------------------------------

//-------------GETTING CURRENT PIXEL COORDINATES-------------
wire [9:0] pix_x;
wire [9:0] pix_y;

pixel_itr show(
	.clk(clk),
   .pix_clk(pix_clk),
	.rst(rst),
	.pix_x(pix_x),
	.pix_y(pix_y),
	.h_sync(h_sync),
	.v_sync(v_sync)
);
//-----------------------------------------------------------

//----------GENERATING WINDOWS LOGO(4 SQUARES)---------------

wire win1, win2, win3, win4;
assign win1 =  (pix_x >= 0 & pix_x <= 71 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 72 & pix_x <= 95 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 96 & pix_x <= 107 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 162 & pix_x <= 215 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 216 & pix_x <= 227 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 252 & pix_x <= 281 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 294 & pix_x <= 305 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 312 & pix_x <= 341 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 342 & pix_x <= 353 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 366 & pix_x <= 377 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 486 & pix_x <= 497 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 72 & pix_x <= 107 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 150 & pix_x <= 185 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 186 & pix_x <= 209 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 210 & pix_x <= 221 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 234 & pix_x <= 263 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 264 & pix_x <= 287 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 288 & pix_x <= 305 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 318 & pix_x <= 335 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 336 & pix_x <= 359 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 480 & pix_x <= 497 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 72 & pix_x <= 119 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 210 & pix_x <= 221 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 240 & pix_x <= 275 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 276 & pix_x <= 305 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 348 & pix_x <= 359 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 486 & pix_x <= 497 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 78 & pix_x <= 101 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 210 & pix_x <= 227 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 228 & pix_x <= 257 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 282 & pix_x <= 299 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 78 & pix_x <= 95 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 156 & pix_x <= 185 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 210 & pix_x <= 233 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 486 & pix_x <= 497 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 78 & pix_x <= 95 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 162 & pix_x <= 185 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 486 & pix_x <= 497 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 78 & pix_x <= 101 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 162 & pix_x <= 179 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 186 & pix_x <= 197 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 78 & pix_x <= 101 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 156 & pix_x <= 173 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 486 & pix_x <= 497 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 78 & pix_x <= 101 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 78 & pix_x <= 95 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 96 & pix_x <= 107 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 108 & pix_x <= 125 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 84 & pix_x <= 113 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 84 & pix_x <= 107 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 84 & pix_x <= 113 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 132 & pix_x <= 149 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 84 & pix_x <= 107 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 108 & pix_x <= 125 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 126 & pix_x <= 143 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 18 & pix_x <= 83 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 84 & pix_x <= 107 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 132 & pix_x <= 143 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 84 & pix_x <= 107 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 90 & pix_x <= 107 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 108 & pix_x <= 131 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 90 & pix_x <= 107 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 108 & pix_x <= 125 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 90 & pix_x <= 113 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 90 & pix_x <= 125 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 150 & pix_x <= 161 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 90 & pix_x <= 113 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 144 & pix_x <= 161 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 96 & pix_x <= 107 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 102 & pix_x <= 113 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 96 & pix_x <= 119 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 126 & pix_x <= 137 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 102 & pix_x <= 125 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 126 & pix_x <= 137 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 30 & pix_x <= 83 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 126 & pix_x <= 137 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 180 & pix_x <= 191 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 132 & pix_x <= 143 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 150 & pix_x <= 161 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 174 & pix_x <= 185 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 78 & pix_x <= 89 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 102 & pix_x <= 113 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 150 & pix_x <= 161 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 36 & pix_x <= 71 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 72 & pix_x <= 83 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 198 & pix_x <= 209 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 54 & pix_x <= 65 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 66 & pix_x <= 77 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 240 & pix_x <= 257 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 324 & pix_x <= 335 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 60 & pix_x <= 71 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 180 & pix_x <= 197 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 186 & pix_x <= 197 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 48 & pix_x <= 65 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 72 & pix_x <= 83 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 132 & pix_x <= 143 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 42 & pix_x <= 59 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 132 & pix_x <= 143 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 42 & pix_x <= 53 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 54 & pix_x <= 65 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 60 & pix_x <= 71 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 42 & pix_x <= 53 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 276 & pix_x <= 293 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 192 & pix_x <= 209 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 222 & pix_x <= 233 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 270 & pix_x <= 293 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 192 & pix_x <= 221 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 270 & pix_x <= 293 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 198 & pix_x <= 227 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 228 & pix_x <= 239 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 264 & pix_x <= 299 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 198 & pix_x <= 233 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 264 & pix_x <= 299 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 192 & pix_x <= 227 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 264 & pix_x <= 299 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 210 & pix_x <= 221 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 264 & pix_x <= 299 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 252 & pix_x <= 305 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 78 & pix_x <= 89 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 246 & pix_x <= 305 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 270 & pix_x <= 293 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 54 & pix_x <= 65 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 54 & pix_x <= 65 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 240 & pix_x <= 263 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 276 & pix_x <= 287 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 252 & pix_x <= 263 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 216 & pix_x <= 227 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 60 & pix_x <= 71 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 264 & pix_x <= 287 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 288 & pix_x <= 299 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 204 & pix_x <= 377 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 198 & pix_x <= 209 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 210 & pix_x <= 239 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 240 & pix_x <= 305 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 306 & pix_x <= 317 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 372 & pix_x <= 383 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 312 & pix_x <= 329 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 378 & pix_x <= 389 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 318 & pix_x <= 329 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 318 & pix_x <= 353 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 192 & pix_x <= 203 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 264 & pix_x <= 275 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 264 & pix_x <= 275 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 174 & pix_x <= 191 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 168 & pix_x <= 197 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 126 & pix_x <= 137 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 168 & pix_x <= 203 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 396 & pix_x <= 407 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 96 & pix_x <= 107 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 168 & pix_x <= 197 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 330 & pix_x <= 341 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 390 & pix_x <= 413 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 78 & pix_x <= 89 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 390 & pix_x <= 401 & pix_y >= 444 & pix_y <= 449);
assign win2 =  (pix_x >= 12 & pix_x <= 29 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 30 & pix_x <= 41 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 78 & pix_x <= 95 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 96 & pix_x <= 185 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 420 & pix_x <= 503 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 510 & pix_x <= 527 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 594 & pix_x <= 599 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 12 & pix_x <= 29 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 30 & pix_x <= 41 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 84 & pix_x <= 95 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 96 & pix_x <= 161 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 246 & pix_x <= 263 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 432 & pix_x <= 509 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 516 & pix_x <= 533 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 12 & pix_x <= 29 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 30 & pix_x <= 41 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 84 & pix_x <= 95 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 96 & pix_x <= 155 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 432 & pix_x <= 503 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 510 & pix_x <= 521 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 12 & pix_x <= 29 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 96 & pix_x <= 149 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 432 & pix_x <= 473 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 480 & pix_x <= 503 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 516 & pix_x <= 527 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 540 & pix_x <= 551 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 24 & pix_x <= 35 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 96 & pix_x <= 143 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 438 & pix_x <= 485 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 540 & pix_x <= 551 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 96 & pix_x <= 143 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 438 & pix_x <= 485 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 102 & pix_x <= 131 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 438 & pix_x <= 455 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 456 & pix_x <= 503 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 540 & pix_x <= 551 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 102 & pix_x <= 143 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 456 & pix_x <= 485 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 102 & pix_x <= 131 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 132 & pix_x <= 143 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 456 & pix_x <= 485 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 540 & pix_x <= 551 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 0 & pix_x <= 11 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 102 & pix_x <= 137 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 462 & pix_x <= 485 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 102 & pix_x <= 137 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 474 & pix_x <= 485 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 102 & pix_x <= 131 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 468 & pix_x <= 485 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 486 & pix_x <= 503 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 558 & pix_x <= 569 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 102 & pix_x <= 137 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 468 & pix_x <= 485 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 504 & pix_x <= 521 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 594 & pix_x <= 599 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 102 & pix_x <= 137 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 456 & pix_x <= 473 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 474 & pix_x <= 485 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 486 & pix_x <= 509 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 594 & pix_x <= 599 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 108 & pix_x <= 137 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 450 & pix_x <= 473 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 474 & pix_x <= 485 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 492 & pix_x <= 515 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 594 & pix_x <= 599 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 450 & pix_x <= 473 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 492 & pix_x <= 515 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 0 & pix_x <= 17 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 108 & pix_x <= 131 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 462 & pix_x <= 473 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 108 & pix_x <= 137 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 462 & pix_x <= 479 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 114 & pix_x <= 149 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 462 & pix_x <= 479 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 114 & pix_x <= 143 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 462 & pix_x <= 479 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 582 & pix_x <= 593 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 0 & pix_x <= 23 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 114 & pix_x <= 143 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 246 & pix_x <= 263 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 462 & pix_x <= 479 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 498 & pix_x <= 509 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 546 & pix_x <= 563 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 114 & pix_x <= 131 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 132 & pix_x <= 149 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 498 & pix_x <= 515 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 114 & pix_x <= 149 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 276 & pix_x <= 287 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 498 & pix_x <= 509 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 114 & pix_x <= 149 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 252 & pix_x <= 263 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 480 & pix_x <= 491 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 498 & pix_x <= 509 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 114 & pix_x <= 149 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 498 & pix_x <= 515 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 120 & pix_x <= 149 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 444 & pix_x <= 467 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 498 & pix_x <= 509 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 120 & pix_x <= 149 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 0 & pix_x <= 29 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 120 & pix_x <= 155 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 450 & pix_x <= 467 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 492 & pix_x <= 515 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 120 & pix_x <= 143 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 228 & pix_x <= 239 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 252 & pix_x <= 263 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 456 & pix_x <= 467 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 582 & pix_x <= 593 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 126 & pix_x <= 155 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 234 & pix_x <= 245 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 252 & pix_x <= 263 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 492 & pix_x <= 509 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 120 & pix_x <= 143 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 240 & pix_x <= 257 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 540 & pix_x <= 551 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 552 & pix_x <= 563 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 120 & pix_x <= 155 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 168 & pix_x <= 185 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 468 & pix_x <= 479 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 126 & pix_x <= 155 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 168 & pix_x <= 185 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 276 & pix_x <= 287 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 552 & pix_x <= 563 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 0 & pix_x <= 35 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 126 & pix_x <= 155 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 468 & pix_x <= 479 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 552 & pix_x <= 563 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 126 & pix_x <= 161 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 450 & pix_x <= 461 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 126 & pix_x <= 161 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 168 & pix_x <= 179 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 468 & pix_x <= 479 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 492 & pix_x <= 503 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 126 & pix_x <= 155 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 168 & pix_x <= 185 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 462 & pix_x <= 479 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 498 & pix_x <= 515 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 546 & pix_x <= 557 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 126 & pix_x <= 167 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 168 & pix_x <= 191 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 540 & pix_x <= 557 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 126 & pix_x <= 167 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 168 & pix_x <= 197 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 132 & pix_x <= 167 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 168 & pix_x <= 197 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 276 & pix_x <= 293 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 132 & pix_x <= 155 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 162 & pix_x <= 209 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 270 & pix_x <= 299 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 438 & pix_x <= 455 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 0 & pix_x <= 41 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 132 & pix_x <= 155 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 162 & pix_x <= 221 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 270 & pix_x <= 299 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 432 & pix_x <= 449 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 450 & pix_x <= 461 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 132 & pix_x <= 155 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 168 & pix_x <= 227 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 264 & pix_x <= 305 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 432 & pix_x <= 449 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 450 & pix_x <= 461 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 132 & pix_x <= 149 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 168 & pix_x <= 251 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 258 & pix_x <= 305 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 342 & pix_x <= 353 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 132 & pix_x <= 161 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 168 & pix_x <= 251 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 252 & pix_x <= 305 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 348 & pix_x <= 371 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 438 & pix_x <= 455 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 132 & pix_x <= 161 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 168 & pix_x <= 185 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 186 & pix_x <= 251 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 252 & pix_x <= 311 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 336 & pix_x <= 365 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 132 & pix_x <= 149 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 174 & pix_x <= 245 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 252 & pix_x <= 305 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 336 & pix_x <= 371 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 414 & pix_x <= 425 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 438 & pix_x <= 455 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 498 & pix_x <= 515 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 0 & pix_x <= 47 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 138 & pix_x <= 161 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 174 & pix_x <= 185 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 186 & pix_x <= 239 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 246 & pix_x <= 323 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 336 & pix_x <= 353 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 432 & pix_x <= 455 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 138 & pix_x <= 155 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 174 & pix_x <= 185 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 186 & pix_x <= 227 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 246 & pix_x <= 323 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 336 & pix_x <= 353 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 138 & pix_x <= 161 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 186 & pix_x <= 197 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 246 & pix_x <= 305 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 312 & pix_x <= 323 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 150 & pix_x <= 167 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 270 & pix_x <= 293 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 306 & pix_x <= 317 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 198 & pix_x <= 209 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 510 & pix_x <= 521 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 180 & pix_x <= 191 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 0 & pix_x <= 53 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 138 & pix_x <= 149 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 276 & pix_x <= 287 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 198 & pix_x <= 209 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 438 & pix_x <= 449 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 162 & pix_x <= 173 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 240 & pix_x <= 257 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 258 & pix_x <= 317 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 0 & pix_x <= 59 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 204 & pix_x <= 377 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 198 & pix_x <= 209 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 216 & pix_x <= 227 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 372 & pix_x <= 383 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 408 & pix_x <= 419 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 444 & pix_x <= 455 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 318 & pix_x <= 347 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 420 & pix_x <= 449 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 450 & pix_x <= 461 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 318 & pix_x <= 347 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 426 & pix_x <= 473 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 192 & pix_x <= 203 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 318 & pix_x <= 353 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 438 & pix_x <= 485 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 180 & pix_x <= 203 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 432 & pix_x <= 503 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 150 & pix_x <= 161 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 168 & pix_x <= 203 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 432 & pix_x <= 521 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 150 & pix_x <= 161 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 162 & pix_x <= 203 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 432 & pix_x <= 539 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 144 & pix_x <= 203 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 432 & pix_x <= 557 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 132 & pix_x <= 203 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 432 & pix_x <= 569 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 114 & pix_x <= 203 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 432 & pix_x <= 593 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 102 & pix_x <= 203 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 396 & pix_x <= 407 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 90 & pix_x <= 203 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 390 & pix_x <= 413 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 78 & pix_x <= 203 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 390 & pix_x <= 413 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 444 & pix_y <= 449);
assign win3 =  (pix_x >= 0 & pix_x <= 203 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 204 & pix_x <= 227 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 252 & pix_x <= 281 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 288 & pix_x <= 305 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 312 & pix_x <= 341 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 342 & pix_x <= 353 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 354 & pix_x <= 389 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 414 & pix_x <= 599 & pix_y >= 0 & pix_y <= 5)| (pix_x >= 0 & pix_x <= 209 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 210 & pix_x <= 227 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 234 & pix_x <= 263 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 264 & pix_x <= 287 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 288 & pix_x <= 305 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 312 & pix_x <= 359 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 366 & pix_x <= 377 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 426 & pix_x <= 599 & pix_y >= 6 & pix_y <= 11)| (pix_x >= 0 & pix_x <= 203 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 204 & pix_x <= 221 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 234 & pix_x <= 305 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 318 & pix_x <= 329 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 330 & pix_x <= 359 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 426 & pix_x <= 599 & pix_y >= 12 & pix_y <= 17)| (pix_x >= 0 & pix_x <= 209 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 210 & pix_x <= 227 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 228 & pix_x <= 263 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 276 & pix_x <= 311 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 330 & pix_x <= 353 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 18 & pix_y <= 23)| (pix_x >= 0 & pix_x <= 185 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 210 & pix_x <= 233 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 294 & pix_x <= 305 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 330 & pix_x <= 341 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 390 & pix_x <= 407 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 24 & pix_y <= 29)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 78 & pix_x <= 185 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 210 & pix_x <= 221 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 222 & pix_x <= 233 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 252 & pix_x <= 263 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 30 & pix_y <= 35)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 78 & pix_x <= 155 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 156 & pix_x <= 179 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 186 & pix_x <= 203 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 216 & pix_x <= 227 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 36 & pix_y <= 41)| (pix_x >= 0 & pix_x <= 101 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 102 & pix_x <= 149 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 156 & pix_x <= 179 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 186 & pix_x <= 197 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 42 & pix_y <= 47)| (pix_x >= 0 & pix_x <= 155 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 174 & pix_x <= 185 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 48 & pix_y <= 53)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 78 & pix_x <= 149 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 54 & pix_y <= 59)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 84 & pix_x <= 149 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 60 & pix_y <= 65)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 78 & pix_x <= 143 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 66 & pix_y <= 71)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 84 & pix_x <= 155 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 156 & pix_x <= 167 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 72 & pix_y <= 77)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 84 & pix_x <= 143 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 78 & pix_y <= 83)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 84 & pix_x <= 107 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 84 & pix_y <= 89)| (pix_x >= 0 & pix_x <= 107 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 90 & pix_y <= 95)| (pix_x >= 0 & pix_x <= 107 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 108 & pix_x <= 143 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 144 & pix_x <= 155 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 96 & pix_y <= 101)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 90 & pix_x <= 149 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 102 & pix_y <= 107)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 90 & pix_x <= 149 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 450 & pix_x <= 599 & pix_y >= 108 & pix_y <= 113)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 90 & pix_x <= 161 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 228 & pix_x <= 269 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 450 & pix_x <= 599 & pix_y >= 114 & pix_y <= 119)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 90 & pix_x <= 161 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 216 & pix_x <= 281 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 450 & pix_x <= 599 & pix_y >= 120 & pix_y <= 125)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 96 & pix_x <= 161 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 210 & pix_x <= 281 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 450 & pix_x <= 599 & pix_y >= 126 & pix_y <= 131)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 114 & pix_x <= 155 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 210 & pix_x <= 293 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 294 & pix_x <= 317 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 324 & pix_x <= 377 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 450 & pix_x <= 599 & pix_y >= 132 & pix_y <= 137)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 114 & pix_x <= 161 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 198 & pix_x <= 383 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 138 & pix_y <= 143)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 96 & pix_x <= 113 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 114 & pix_x <= 161 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 192 & pix_x <= 389 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 144 & pix_y <= 149)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 96 & pix_x <= 155 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 186 & pix_x <= 395 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 150 & pix_y <= 155)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 96 & pix_x <= 155 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 186 & pix_x <= 395 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 156 & pix_y <= 161)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 96 & pix_x <= 155 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 186 & pix_x <= 389 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 162 & pix_y <= 167)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 96 & pix_x <= 119 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 120 & pix_x <= 155 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 180 & pix_x <= 389 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 168 & pix_y <= 173)| (pix_x >= 0 & pix_x <= 95 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 120 & pix_x <= 155 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 180 & pix_x <= 395 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 174 & pix_y <= 179)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 102 & pix_x <= 119 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 120 & pix_x <= 161 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 174 & pix_x <= 395 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 180 & pix_y <= 185)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 120 & pix_x <= 155 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 168 & pix_x <= 407 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 186 & pix_y <= 191)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 102 & pix_x <= 161 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 168 & pix_x <= 419 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 444 & pix_x <= 599 & pix_y >= 192 & pix_y <= 197)| (pix_x >= 0 & pix_x <= 95 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 102 & pix_x <= 161 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 168 & pix_x <= 419 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 198 & pix_y <= 203)| (pix_x >= 0 & pix_x <= 95 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 102 & pix_x <= 161 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 168 & pix_x <= 203 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 204 & pix_x <= 221 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 228 & pix_x <= 401 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 402 & pix_x <= 413 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 426 & pix_x <= 599 & pix_y >= 204 & pix_y <= 209)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 84 & pix_x <= 95 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 108 & pix_x <= 119 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 126 & pix_x <= 161 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 168 & pix_x <= 191 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 258 & pix_x <= 311 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 396 & pix_x <= 419 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 210 & pix_y <= 215)| (pix_x >= 0 & pix_x <= 95 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 108 & pix_x <= 125 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 126 & pix_x <= 161 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 168 & pix_x <= 203 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 264 & pix_x <= 305 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 396 & pix_x <= 413 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 216 & pix_y <= 221)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 108 & pix_x <= 125 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 126 & pix_x <= 167 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 168 & pix_x <= 233 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 264 & pix_x <= 299 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 378 & pix_x <= 395 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 396 & pix_x <= 419 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 222 & pix_y <= 227)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 126 & pix_x <= 215 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 216 & pix_x <= 227 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 270 & pix_x <= 299 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 354 & pix_x <= 365 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 384 & pix_x <= 419 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 228 & pix_y <= 233)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 66 & pix_x <= 77 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 78 & pix_x <= 89 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 108 & pix_x <= 203 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 264 & pix_x <= 305 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 342 & pix_x <= 353 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 378 & pix_x <= 413 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 426 & pix_x <= 599 & pix_y >= 234 & pix_y <= 239)| (pix_x >= 0 & pix_x <= 65 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 66 & pix_x <= 77 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 108 & pix_x <= 203 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 264 & pix_x <= 305 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 384 & pix_x <= 419 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 420 & pix_x <= 431 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 240 & pix_y <= 245)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 72 & pix_x <= 89 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 114 & pix_x <= 215 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 264 & pix_x <= 305 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 378 & pix_x <= 419 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 420 & pix_x <= 599 & pix_y >= 246 & pix_y <= 251)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 114 & pix_x <= 125 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 132 & pix_x <= 221 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 222 & pix_x <= 233 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 240 & pix_x <= 305 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 366 & pix_x <= 413 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 414 & pix_x <= 599 & pix_y >= 252 & pix_y <= 257)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 72 & pix_x <= 83 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 84 & pix_x <= 95 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 132 & pix_x <= 335 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 348 & pix_x <= 359 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 360 & pix_x <= 419 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 420 & pix_x <= 599 & pix_y >= 258 & pix_y <= 263)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 132 & pix_x <= 413 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 414 & pix_x <= 599 & pix_y >= 264 & pix_y <= 269)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 120 & pix_x <= 131 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 132 & pix_x <= 413 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 414 & pix_x <= 599 & pix_y >= 270 & pix_y <= 275)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 132 & pix_x <= 407 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 408 & pix_x <= 599 & pix_y >= 276 & pix_y <= 281)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 132 & pix_x <= 407 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 408 & pix_x <= 599 & pix_y >= 282 & pix_y <= 287)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 78 & pix_x <= 89 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 132 & pix_x <= 407 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 408 & pix_x <= 599 & pix_y >= 288 & pix_y <= 293)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 132 & pix_x <= 401 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 294 & pix_y <= 299)| (pix_x >= 0 & pix_x <= 83 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 138 & pix_x <= 395 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 300 & pix_y <= 305)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 138 & pix_x <= 395 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 306 & pix_y <= 311)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 126 & pix_x <= 137 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 138 & pix_x <= 389 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 312 & pix_y <= 317)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 138 & pix_x <= 263 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 270 & pix_x <= 299 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 312 & pix_x <= 389 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 318 & pix_y <= 323)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 138 & pix_x <= 233 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 234 & pix_x <= 263 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 270 & pix_x <= 293 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 318 & pix_x <= 389 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 396 & pix_x <= 599 & pix_y >= 324 & pix_y <= 329)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 138 & pix_x <= 227 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 240 & pix_x <= 275 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 276 & pix_x <= 293 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 348 & pix_x <= 383 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 384 & pix_x <= 395 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 396 & pix_x <= 599 & pix_y >= 330 & pix_y <= 335)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 144 & pix_x <= 227 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 240 & pix_x <= 293 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 354 & pix_x <= 371 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 384 & pix_x <= 395 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 396 & pix_x <= 599 & pix_y >= 336 & pix_y <= 341)| (pix_x >= 0 & pix_x <= 89 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 144 & pix_x <= 227 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 258 & pix_x <= 305 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 306 & pix_x <= 317 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 354 & pix_x <= 389 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 390 & pix_x <= 599 & pix_y >= 342 & pix_y <= 347)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 144 & pix_x <= 233 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 234 & pix_x <= 251 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 264 & pix_x <= 281 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 282 & pix_x <= 299 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 354 & pix_x <= 371 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 378 & pix_x <= 389 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 390 & pix_x <= 599 & pix_y >= 348 & pix_y <= 353)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 144 & pix_x <= 269 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 306 & pix_x <= 341 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 342 & pix_x <= 365 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 390 & pix_x <= 599 & pix_y >= 354 & pix_y <= 359)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 144 & pix_x <= 359 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 390 & pix_x <= 599 & pix_y >= 360 & pix_y <= 365)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 144 & pix_x <= 377 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 378 & pix_x <= 389 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 396 & pix_x <= 599 & pix_y >= 366 & pix_y <= 371)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 144 & pix_x <= 317 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 372 & pix_x <= 389 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 402 & pix_x <= 599 & pix_y >= 372 & pix_y <= 377)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 312 & pix_x <= 347 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 378 & pix_x <= 389 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 414 & pix_x <= 599 & pix_y >= 378 & pix_y <= 383)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 240 & pix_x <= 251 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 312 & pix_x <= 347 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 348 & pix_x <= 359 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 360 & pix_x <= 371 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 426 & pix_x <= 599 & pix_y >= 384 & pix_y <= 389)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 246 & pix_x <= 257 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 318 & pix_x <= 365 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 438 & pix_x <= 599 & pix_y >= 390 & pix_y <= 395)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 396 & pix_y <= 401)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 258 & pix_x <= 269 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 402 & pix_y <= 407)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 258 & pix_x <= 275 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 408 & pix_y <= 413)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 150 & pix_x <= 203 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 258 & pix_x <= 275 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 414 & pix_y <= 419)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 132 & pix_x <= 203 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 264 & pix_x <= 281 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 420 & pix_y <= 425)| (pix_x >= 0 & pix_x <= 71 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 114 & pix_x <= 203 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 270 & pix_x <= 281 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 426 & pix_y <= 431)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 108 & pix_x <= 203 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 396 & pix_x <= 407 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 432 & pix_y <= 437)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 90 & pix_x <= 203 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 330 & pix_x <= 341 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 390 & pix_x <= 413 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 438 & pix_y <= 443)| (pix_x >= 0 & pix_x <= 77 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 78 & pix_x <= 203 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 336 & pix_x <= 347 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 384 & pix_x <= 413 & pix_y >= 444 & pix_y <= 449)| (pix_x >= 432 & pix_x <= 599 & pix_y >= 444 & pix_y <= 449);

//assign win1 = (pix_y > 400) & (pix_y < 450);
//assign win2 = (pix_x > 620) & (pix_x < 630);
//assign win3 = (pix_x > 20) & (pix_x< 640); 
//becomes a 853x480 display on 16:9

assign r_out = win1;
assign g_out = win2;
assign b_out = win3;
//assign temp = win4;

//-----------------------------------------------------------


endmodule
