VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  CAPACITANCE PICOFARADS 1 ;
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
LAYER Oxide
  TYPE MASTERSLICE ;
END Oxide

LAYER Poly
  TYPE MASTERSLICE ;
END Poly

LAYER Nhvt
  TYPE IMPLANT ;
END Nhvt

LAYER Nimp
  TYPE IMPLANT ;
  WIDTH 0.24 ;
  SPACING 0.24 ;
END Nimp

LAYER Phvt
  TYPE IMPLANT ;
END Phvt

LAYER Pimp
  TYPE IMPLANT ;
  WIDTH 0.24 ;
  SPACING 0.24 ;
  SPACING 0 LAYER Nimp ;
END Pimp

LAYER Nzvt
  TYPE IMPLANT ;
  WIDTH 0.7 ;
  SPACING 0.6 ;
END Nzvt

LAYER SiProt
  TYPE IMPLANT ;
  WIDTH 0.44 ;
  SPACING 0.44 ;
END SiProt

LAYER Cont
  TYPE CUT ;
  SPACING 0.14 ;
  SPACING 0.16 ADJACENTCUTS 3 WITHIN 0.17 ;
  WIDTH 0.12 ;
  ENCLOSURE BELOW 0.04 0.06 ;
  ENCLOSURE ABOVE 0 0.06 ;
  ANTENNAMODEL OXIDE1 ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.12 ;
  AREA 0.07 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.12 0.12 0.12 0.12 0.12 0.12 
    WIDTH 0.18 0.12 0.18 0.18 0.18 0.18 0.18 
    WIDTH 1.5 0.18 0.18 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.12 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 1 WIDTH 0.14 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.08 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.3 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal1

LAYER Via1
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal2

LAYER Via2
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal3

LAYER Via3
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal4

LAYER Via4
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 ;
  MINIMUMCUT 2 WIDTH 0.4 ;
  MINIMUMCUT 4 WIDTH 1 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal5

LAYER Via5
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 ;
  MINIMUMCUT 2 WIDTH 0.4 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 1 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.6 FROMABOVE ;
  MINIMUMCUT 4 WIDTH 4 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal6

LAYER Via6
  TYPE CUT ;
  SPACING 0.15 ;
  SPACING 0.2 ADJACENTCUTS 3 WITHIN 0.21 ;
  WIDTH 0.14 ;
  ENCLOSURE BELOW 0.005 0.06 ;
  ENCLOSURE ABOVE 0.005 0.06 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.1 ;
END Via6

LAYER Metal7
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.29 0.29 ;
  WIDTH 0.14 ;
  AREA 0.08 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 0.5585 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.14 0.14 0.14 0.14 0.14 0.14 
    WIDTH 0.2 0.14 0.2 0.2 0.2 0.2 0.2 
    WIDTH 1.5 0.2 0.2 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 1 WIDTH 0.14 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.6 FROMBELOW ;
  MINIMUMCUT 4 WIDTH 4 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.06 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 0.36 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 2 ;
END Metal7

LAYER Via7
  TYPE CUT ;
  SPACING 0.36 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.55 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.03 0.08 ;
  ENCLOSURE ABOVE 0.05 0.1 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.8 ;
END Via7

LAYER Metal8
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.87 0.87 ;
  WIDTH 0.44 ;
  AREA 0.2 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.4 0.4 0.4 0.4 0.4 
    WIDTH 1.5 0.4 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MINIMUMCUT 2 WIDTH 2 FROMABOVE LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.02 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 8 ;
END Metal8

LAYER Via8
  TYPE CUT ;
  SPACING 0.36 ;
  SPACING 0.54 ADJACENTCUTS 3 WITHIN 0.55 ;
  WIDTH 0.36 ;
  ENCLOSURE BELOW 0.03 0.08 ;
  ENCLOSURE ABOVE 0.05 0.1 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 25 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 25 ) ( 0.099 25 ) ( 0.1 1025 ) ( 1 1250 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.8 ;
END Via8

LAYER Metal9
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.87 0.87 ;
  WIDTH 0.44 ;
  AREA 0.2 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.4985 2.9985 4.4985 7.4985 
    WIDTH 0 0.4 0.4 0.4 0.4 0.4 
    WIDTH 1.5 0.4 0.5 0.5 0.5 0.5 
    WIDTH 3 0.5 0.5 0.9 0.9 0.9 
    WIDTH 4.5 0.9 0.9 0.9 1.5 1.5 
    WIDTH 7.5 1.5 1.5 1.5 1.5 2.5 ;
  MINIMUMCUT 2 WIDTH 2 FROMBELOW LENGTH 20 WITHIN 5 ;
  MAXWIDTH 12 ;
  RESISTANCE RPERSQ 0.02 ;
  CAPACITANCE CPERSQDIST 0.0002 ;
  THICKNESS 1 ;
  EDGECAPACITANCE 0.0002 ;
  MINIMUMDENSITY 20 ;
  MAXIMUMDENSITY 65 ;
  DENSITYCHECKWINDOW 120 120 ;
  DENSITYCHECKSTEP 60 ;
  ANTENNAMODEL OXIDE1 ;
    ANTENNAAREARATIO 475 ;
    ANTENNACUMAREARATIO 1200 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1200 ) ( 0.099 1200 ) ( 0.1 55750 ) ( 1 62500 ) ) ;
  DCCURRENTDENSITY AVERAGE 8 ;
END Metal9

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

MAXVIASTACK 4 RANGE Metal1 Metal7 ;
VIA VIA1X DEFAULT
  LAYER Metal1 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA1X

VIA VIA1V DEFAULT
  LAYER Metal1 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA1V

VIA VIA1H DEFAULT
  LAYER Metal1 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA1H

VIA VIA1XR90 DEFAULT
  LAYER Metal1 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA1XR90

VIA VIA1_2CUT_E DEFAULT
  LAYER Metal1 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_E

VIA VIA1_2CUT_W DEFAULT
  LAYER Metal1 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via1 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_W

VIA VIA1_2CUT_N DEFAULT
  LAYER Metal1 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_N

VIA VIA1_2CUT_S DEFAULT
  LAYER Metal1 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via1 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal2 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_S

VIA VIA1_2X2CUT DEFAULT
  LAYER Metal1 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  LAYER Via1 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal2 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  RESISTANCE 0.35 ;
END VIA1_2X2CUT

VIA VIA2X DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA2X

VIA VIA2H DEFAULT
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA2H

VIA VIA2V DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA2V

VIA VIA2XR90 DEFAULT
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA2XR90

VIA VIA2TOS DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA2TOS

VIA VIA2TOS_S DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA2TOS_S

VIA VIA2TOS_N DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA2TOS_N

VIA VIA2_2CUT_N DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_N

VIA VIA2_2CUT_S DEFAULT
  LAYER Metal2 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via2 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_S

VIA VIA2_2CUT_E DEFAULT
  LAYER Metal2 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_E

VIA VIA2_2CUT_W DEFAULT
  LAYER Metal2 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via2 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal3 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_W

VIA VIA2_2X2CUT DEFAULT
  LAYER Metal2 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  LAYER Via2 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal3 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  RESISTANCE 0.35 ;
END VIA2_2X2CUT

VIA VIA3X DEFAULT
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA3X

VIA VIA3H DEFAULT
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA3H

VIA VIA3V DEFAULT
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA3V

VIA VIA3XR90 DEFAULT
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA3XR90

VIA VIA3TOS_E DEFAULT
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.41 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA3TOS_E

VIA VIA3TOS_W DEFAULT
  LAYER Metal3 ;
    RECT -0.41 -0.075 0.13 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA3TOS_W

VIA VIA3TOS DEFAULT
  LAYER Metal3 ;
    RECT -0.27 -0.075 0.27 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA3TOS

VIA VIA3_2CUT_E DEFAULT
  LAYER Metal3 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_E

VIA VIA3_2CUT_W DEFAULT
  LAYER Metal3 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via3 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_W

VIA VIA3_2CUT_N DEFAULT
  LAYER Metal3 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_N

VIA VIA3_2CUT_S DEFAULT
  LAYER Metal3 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via3 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal4 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_S

VIA VIA3_2X2CUT DEFAULT
  LAYER Metal3 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  LAYER Via3 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal4 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  RESISTANCE 0.35 ;
END VIA3_2X2CUT

VIA VIA4X DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA4X

VIA VIA4H DEFAULT
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA4H

VIA VIA4V DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA4V

VIA VIA4XR90 DEFAULT
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA4XR90

VIA VIA4TOS DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA4TOS

VIA VIA4TOS_S DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA4TOS_S

VIA VIA4TOS_N DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA4TOS_N

VIA VIA4_2CUT_N DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_N

VIA VIA4_2CUT_S DEFAULT
  LAYER Metal4 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via4 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_S

VIA VIA4_2CUT_E DEFAULT
  LAYER Metal4 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_E

VIA VIA4_2CUT_W DEFAULT
  LAYER Metal4 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via4 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal5 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_W

VIA VIA4_2X2CUT DEFAULT
  LAYER Metal4 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  LAYER Via4 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal5 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  RESISTANCE 0.35 ;
END VIA4_2X2CUT

VIA VIA5X DEFAULT
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA5X

VIA VIA5H DEFAULT
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA5H

VIA VIA5V DEFAULT
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA5V

VIA VIA5XR90 DEFAULT
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA5XR90

VIA VIA5TOS_E DEFAULT
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.41 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA5TOS_E

VIA VIA5TOS_W DEFAULT
  LAYER Metal5 ;
    RECT -0.41 -0.075 0.13 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA5TOS_W

VIA VIA5TOS DEFAULT
  LAYER Metal5 ;
    RECT -0.27 -0.075 0.27 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA5TOS

VIA VIA5_2CUT_E DEFAULT
  LAYER Metal5 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_E

VIA VIA5_2CUT_W DEFAULT
  LAYER Metal5 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via5 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_W

VIA VIA5_2CUT_N DEFAULT
  LAYER Metal5 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_N

VIA VIA5_2CUT_S DEFAULT
  LAYER Metal5 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via5 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal6 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_S

VIA VIA5_2X2CUT DEFAULT
  LAYER Metal5 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  LAYER Via5 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal6 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  RESISTANCE 0.35 ;
END VIA5_2X2CUT

VIA VIA6X DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA6X

VIA VIA6H DEFAULT
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA6H

VIA VIA6V DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA6V

VIA VIA6XR90 DEFAULT
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.075 -0.13 0.075 0.13 ;
  RESISTANCE 1.4 ;
END VIA6XR90

VIA VIA6TOS DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.27 0.075 0.27 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA6TOS

VIA VIA6TOS_S DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.41 0.075 0.13 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA6TOS_S

VIA VIA6TOS_N DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.41 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.13 0.075 ;
  RESISTANCE 1.4 ;
END VIA6TOS_N

VIA VIA6_2CUT_N DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT -0.07 0.22 0.07 0.36 ;
  LAYER Metal7 ;
    RECT -0.075 -0.13 0.075 0.42 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_N

VIA VIA6_2CUT_S DEFAULT
  LAYER Metal6 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  LAYER Via6 ;
    RECT -0.07 -0.36 0.07 -0.22 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.075 -0.42 0.075 0.13 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_S

VIA VIA6_2CUT_E DEFAULT
  LAYER Metal6 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    RECT 0.22 -0.07 0.36 0.07 ;
  LAYER Metal7 ;
    RECT -0.13 -0.075 0.42 0.075 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_E

VIA VIA6_2CUT_W DEFAULT
  LAYER Metal6 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  LAYER Via6 ;
    RECT -0.36 -0.07 -0.22 0.07 ;
    RECT -0.07 -0.07 0.07 0.07 ;
  LAYER Metal7 ;
    RECT -0.42 -0.075 0.13 0.075 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_W

VIA VIA6_2X2CUT DEFAULT
  LAYER Metal6 ;
    RECT -0.22 -0.275 0.22 0.275 ;
  LAYER Via6 ;
    RECT 0.075 0.075 0.215 0.215 ;
    RECT -0.215 0.075 -0.075 0.215 ;
    RECT -0.215 -0.215 -0.075 -0.075 ;
    RECT 0.075 -0.215 0.215 -0.075 ;
  LAYER Metal7 ;
    RECT -0.275 -0.22 0.275 0.22 ;
  RESISTANCE 0.35 ;
END VIA6_2X2CUT

VIA VIA7X DEFAULT
  LAYER Metal7 ;
    RECT -0.26 -0.21 0.26 0.21 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -0.23 -0.28 0.23 0.28 ;
  RESISTANCE 0.35 ;
END VIA7X

VIA VIA7V DEFAULT
  LAYER Metal7 ;
    RECT -0.21 -0.26 0.21 0.26 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -0.23 -0.28 0.23 0.28 ;
  RESISTANCE 0.35 ;
END VIA7V

VIA VIA7H DEFAULT
  LAYER Metal7 ;
    RECT -0.26 -0.21 0.26 0.21 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -0.28 -0.23 0.28 0.23 ;
  RESISTANCE 0.35 ;
END VIA7H

VIA VIA7XR90 DEFAULT
  LAYER Metal7 ;
    RECT -0.21 -0.26 0.21 0.26 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -0.23 -0.28 0.23 0.28 ;
  RESISTANCE 0.35 ;
END VIA7XR90

VIA VIA7_2CUT_E DEFAULT
  LAYER Metal7 ;
    RECT -0.26 -0.21 0.98 0.21 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    RECT 0.54 -0.18 0.9 0.18 ;
  LAYER Metal8 ;
    RECT -0.28 -0.23 1 0.23 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_E

VIA VIA7_2CUT_W DEFAULT
  LAYER Metal7 ;
    RECT -0.98 -0.21 0.26 0.21 ;
  LAYER Via7 ;
    RECT -0.9 -0.18 -0.54 0.18 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -1 -0.23 0.28 0.23 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_W

VIA VIA7_2CUT_N DEFAULT
  LAYER Metal7 ;
    RECT -0.21 -0.26 0.21 0.98 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    RECT -0.18 0.54 0.18 0.9 ;
  LAYER Metal8 ;
    RECT -0.23 -0.28 0.23 1 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_N

VIA VIA7_2CUT_S DEFAULT
  LAYER Metal7 ;
    RECT -0.21 -0.98 0.21 0.26 ;
  LAYER Via7 ;
    RECT -0.18 -0.9 0.18 -0.54 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal8 ;
    RECT -0.23 -1 0.23 0.28 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_S

VIA VIA7_2X2CUT DEFAULT
  LAYER Metal7 ;
    RECT -0.71 -0.66 0.71 0.66 ;
  LAYER Via7 ;
    RECT 0.27 0.27 0.63 0.63 ;
    RECT -0.63 0.27 -0.27 0.63 ;
    RECT -0.63 -0.63 -0.27 -0.27 ;
    RECT 0.27 -0.63 0.63 -0.27 ;
  LAYER Metal8 ;
    RECT -0.68 -0.73 0.68 0.73 ;
  RESISTANCE 0.0875 ;
END VIA7_2X2CUT

VIA VIA8X DEFAULT
  LAYER Metal8 ;
    RECT -0.23 -0.26 0.23 0.26 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -0.28 -0.23 0.28 0.23 ;
  RESISTANCE 0.35 ;
END VIA8X

VIA VIA8H DEFAULT
  LAYER Metal8 ;
    RECT -0.26 -0.23 0.26 0.23 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -0.28 -0.23 0.28 0.23 ;
  RESISTANCE 0.35 ;
END VIA8H

VIA VIA8V DEFAULT
  LAYER Metal8 ;
    RECT -0.23 -0.26 0.23 0.26 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -0.23 -0.28 0.23 0.28 ;
  RESISTANCE 0.35 ;
END VIA8V

VIA VIA8XR90 DEFAULT
  LAYER Metal8 ;
    RECT -0.26 -0.23 0.26 0.23 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -0.23 -0.28 0.23 0.28 ;
  RESISTANCE 0.35 ;
END VIA8XR90

VIA VIA8_2CUT_E DEFAULT
  LAYER Metal8 ;
    RECT -0.26 -0.23 0.98 0.23 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    RECT 0.54 -0.18 0.9 0.18 ;
  LAYER Metal9 ;
    RECT -0.28 -0.23 1 0.23 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_E

VIA VIA8_2CUT_W DEFAULT
  LAYER Metal8 ;
    RECT -0.98 -0.23 0.26 0.23 ;
  LAYER Via8 ;
    RECT -0.9 -0.18 -0.54 0.18 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -1 -0.23 0.28 0.23 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_W

VIA VIA8_2CUT_N DEFAULT
  LAYER Metal8 ;
    RECT -0.23 -0.26 0.23 0.98 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    RECT -0.18 0.54 0.18 0.9 ;
  LAYER Metal9 ;
    RECT -0.23 -0.28 0.23 1 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_N

VIA VIA8_2CUT_S DEFAULT
  LAYER Metal8 ;
    RECT -0.23 -0.98 0.23 0.26 ;
  LAYER Via8 ;
    RECT -0.18 -0.9 0.18 -0.54 ;
    RECT -0.18 -0.18 0.18 0.18 ;
  LAYER Metal9 ;
    RECT -0.23 -1 0.23 0.28 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_S

VIA VIA8_2X2CUT DEFAULT
  LAYER Metal8 ;
    RECT -0.66 -0.71 0.66 0.71 ;
  LAYER Via8 ;
    RECT 0.27 0.27 0.63 0.63 ;
    RECT -0.63 0.27 -0.27 0.63 ;
    RECT -0.63 -0.63 -0.27 -0.27 ;
    RECT 0.27 -0.63 0.63 -0.27 ;
  LAYER Metal9 ;
    RECT -0.73 -0.68 0.73 0.68 ;
  RESISTANCE 0.0875 ;
END VIA8_2X2CUT

VIA VIA1_2CUT_H
  LAYER Metal1 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via1 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal2 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_H

VIA VIA1_2CUT_V
  LAYER Metal1 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via1 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal2 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA1_2CUT_V

VIA VIA2_2CUT_H
  LAYER Metal2 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via2 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal3 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_H

VIA VIA2_2CUT_V
  LAYER Metal2 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via2 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal3 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA2_2CUT_V

VIA VIA3_2CUT_H
  LAYER Metal3 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via3 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal4 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_H

VIA VIA3_2CUT_V
  LAYER Metal3 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via3 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal4 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA3_2CUT_V

VIA VIA4_2CUT_H
  LAYER Metal4 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via4 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal5 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_H

VIA VIA4_2CUT_V
  LAYER Metal4 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via4 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal5 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA4_2CUT_V

VIA VIA5_2CUT_H
  LAYER Metal5 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via5 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal6 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_H

VIA VIA5_2CUT_V
  LAYER Metal5 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via5 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal6 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA5_2CUT_V

VIA VIA6_2CUT_H
  LAYER Metal6 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  LAYER Via6 ;
    RECT -0.215 -0.07 -0.075 0.07 ;
    RECT 0.075 -0.07 0.215 0.07 ;
  LAYER Metal7 ;
    RECT -0.275 -0.075 0.275 0.075 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_H

VIA VIA6_2CUT_V
  LAYER Metal6 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  LAYER Via6 ;
    RECT -0.07 -0.215 0.07 -0.075 ;
    RECT -0.07 0.075 0.07 0.215 ;
  LAYER Metal7 ;
    RECT -0.075 -0.275 0.075 0.275 ;
  RESISTANCE 0.7 ;
END VIA6_2CUT_V

VIA VIA7_2CUT_H
  LAYER Metal7 ;
    RECT -0.62 -0.21 0.62 0.21 ;
  LAYER Via7 ;
    RECT -0.54 -0.18 -0.18 0.18 ;
    RECT 0.18 -0.18 0.54 0.18 ;
  LAYER Metal8 ;
    RECT -0.64 -0.23 0.64 0.23 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_H

VIA VIA7_2CUT_V
  LAYER Metal7 ;
    RECT -0.21 -0.62 0.21 0.62 ;
  LAYER Via7 ;
    RECT -0.18 -0.54 0.18 -0.18 ;
    RECT -0.18 0.18 0.18 0.54 ;
  LAYER Metal8 ;
    RECT -0.23 -0.64 0.23 0.64 ;
  RESISTANCE 0.175 ;
END VIA7_2CUT_V

VIA VIA8_2CUT_H
  LAYER Metal8 ;
    RECT -0.62 -0.23 0.62 0.23 ;
  LAYER Via8 ;
    RECT -0.54 -0.18 -0.18 0.18 ;
    RECT 0.18 -0.18 0.54 0.18 ;
  LAYER Metal9 ;
    RECT -0.64 -0.23 0.64 0.23 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_H

VIA VIA8_2CUT_V
  LAYER Metal8 ;
    RECT -0.23 -0.62 0.23 0.62 ;
  LAYER Via8 ;
    RECT -0.18 -0.54 0.18 -0.18 ;
    RECT -0.18 0.18 0.18 0.54 ;
  LAYER Metal9 ;
    RECT -0.23 -0.64 0.23 0.64 ;
  RESISTANCE 0.175 ;
END VIA8_2CUT_V

VIARULE VIA1ARRAY GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA1ARRAY

VIARULE VIA2ARRAY GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA2ARRAY

VIARULE VIA3ARRAY GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA3ARRAY

VIARULE VIA4ARRAY GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA4ARRAY

VIARULE VIA5ARRAY GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA5ARRAY

VIARULE VIA6ARRAY GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.06 0.005 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
    RESISTANCE 1.400000 ;
END VIA6ARRAY

VIARULE VIA7ARRAY GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.08 0.03 ;
  LAYER Metal8 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.9 BY 0.9 ;
    RESISTANCE 0.350000 ;
END VIA7ARRAY

VIARULE VIA8ARRAY GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.04 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.1 0.05 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.9 BY 0.9 ;
    RESISTANCE 0.350000 ;
END VIA8ARRAY

VIARULE M9_M8v GENERATE DEFAULT
  LAYER Metal8 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8v

VIARULE M8_M7v GENERATE DEFAULT
  LAYER Metal7 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7v

VIARULE M7_M6v GENERATE DEFAULT
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M7_M6v

VIARULE M6_M5v GENERATE DEFAULT
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M6_M5v

VIARULE M5_M4v GENERATE DEFAULT
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M5_M4v

VIARULE M4_M3v GENERATE DEFAULT
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M4_M3v

VIARULE M3_M2v GENERATE DEFAULT
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M3_M2v

VIARULE M2_M1v GENERATE DEFAULT
  LAYER Metal1 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.29 BY 0.29 ;
END M2_M1v

VIARULE M1_POv GENERATE DEFAULT
  LAYER Poly ;
    ENCLOSURE 0.04 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.26 BY 0.26 ;
END M1_POv

VIARULE M1_DIFF GENERATE DEFAULT
  LAYER Oxide ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_DIFF

VIARULE M1_PSUB GENERATE DEFAULT
  LAYER Oxide ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_PSUB

VIARULE M1_PIMP GENERATE DEFAULT
  LAYER Oxide ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_PIMP

VIARULE M1_NIMP GENERATE DEFAULT
  LAYER Oxide ;
    ENCLOSURE 0.07 0.07 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_NIMP

VIARULE M1_NWELL GENERATE DEFAULT
  LAYER Oxide ;
    ENCLOSURE 0.07 0.07 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_NWELL

VIARULE M9_M8 GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8

VIARULE M8_M7 GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.08 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7

VIARULE M7_M6 GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M7_M6

VIARULE M6_M5 GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M6_M5

VIARULE M5_M4 GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M5_M4

VIARULE M4_M3 GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M4_M3

VIARULE M3_M2 GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M2_M1

VIARULE M1_PO GENERATE
  LAYER Poly ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0.06 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_PO

VIARULE M9_M8c GENERATE
  LAYER Metal8 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal9 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via8 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M9_M8c

VIARULE M8_M7c GENERATE
  LAYER Metal7 ;
    ENCLOSURE 0.03 0.08 ;
  LAYER Metal8 ;
    ENCLOSURE 0.05 0.1 ;
  LAYER Via7 ;
    RECT -0.18 -0.18 0.18 0.18 ;
    SPACING 0.72 BY 0.72 ;
END M8_M7c

VIARULE M7_M6c GENERATE
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal7 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via6 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M7_M6c

VIARULE M6_M5c GENERATE
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal6 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via5 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M6_M5c

VIARULE M5_M4c GENERATE
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal5 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via4 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M5_M4c

VIARULE M4_M3c GENERATE
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal4 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via3 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M4_M3c

VIARULE M3_M2c GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal3 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via2 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M3_M2c

VIARULE M2_M1c GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Metal2 ;
    ENCLOSURE 0.005 0.06 ;
  LAYER Via1 ;
    RECT -0.07 -0.07 0.07 0.07 ;
    SPACING 0.34 BY 0.34 ;
END M2_M1c

VIARULE M1_DIFFc GENERATE
  LAYER Oxide ;
    ENCLOSURE 0.1 0.1 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_DIFFc

VIARULE M1_POLYc GENERATE
  LAYER Poly ;
    ENCLOSURE 0.04 0.06 ;
  LAYER Metal1 ;
    ENCLOSURE 0 0.06 ;
  LAYER Cont ;
    RECT -0.06 -0.06 0.06 0.06 ;
    SPACING 0.28 BY 0.28 ;
END M1_POLYc

SPACING
  SAMENET Oxide Oxide 0.15 ;
  SAMENET Poly Poly 0.12 ;
  SAMENET Cont Cont 0.14 ;
  SAMENET Metal1 Metal1 0.12 ;
  SAMENET Via1 Via1 0.15 ;
  SAMENET Metal2 Metal2 0.14 ;
  SAMENET Via2 Via2 0.15 ;
  SAMENET Metal3 Metal3 0.14 ;
  SAMENET Via3 Via3 0.15 ;
  SAMENET Metal4 Metal4 0.14 ;
  SAMENET Via4 Via4 0.15 ;
  SAMENET Metal5 Metal5 0.14 ;
  SAMENET Via5 Via5 0.15 ;
  SAMENET Metal6 Metal6 0.14 ;
  SAMENET Via6 Via6 0.15 ;
  SAMENET Metal7 Metal7 0.14 ;
  SAMENET Via7 Via7 0.36 ;
  SAMENET Metal8 Metal8 0.4 ;
  SAMENET Via8 Via8 0.36 ;
  SAMENET Metal9 Metal9 0.4 ;
END SPACING

NONDEFAULTRULE LEFDefaultRouteSpec_gpdk090
  LAYER Metal1
    WIDTH 0.12 ;
  END Metal1
  LAYER Metal2
    WIDTH 0.14 ;
  END Metal2
  LAYER Metal3
    WIDTH 0.14 ;
  END Metal3
  LAYER Metal4
    WIDTH 0.14 ;
  END Metal4
  LAYER Metal5
    WIDTH 0.14 ;
  END Metal5
  LAYER Metal6
    WIDTH 0.14 ;
  END Metal6
  LAYER Metal7
    WIDTH 0.14 ;
  END Metal7
  LAYER Metal8
    WIDTH 0.44 ;
  END Metal8
  LAYER Metal9
    WIDTH 0.44 ;
  END Metal9
  USEVIARULE M1_POv ;
  USEVIARULE M2_M1v ;
  USEVIARULE M3_M2v ;
  USEVIARULE M4_M3v ;
  USEVIARULE M5_M4v ;
  USEVIARULE M6_M5v ;
  USEVIARULE M7_M6v ;
  USEVIARULE M8_M7v ;
  USEVIARULE M9_M8v ;
  USEVIARULE M1_NWELL ;
  USEVIARULE M1_PSUB ;
  USEVIARULE M1_NIMP ;
  USEVIARULE M1_PIMP ;
  USEVIARULE M1_DIFF ;
END LEFDefaultRouteSpec_gpdk090
SITE corner
  CLASS PAD ;
  SYMMETRY X Y R90 ;
  SIZE 160 BY 160 ;
END corner

SITE gsclib090site
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.29 BY 2.61 ;
END gsclib090site

SITE pad
  CLASS PAD ;
  SYMMETRY X Y R90 ;
  SIZE 0.005 BY 160 ;
END pad

MACRO OAI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X4 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.795 1.075 3.375 1.195 ;
        RECT 0.68 1.04 2.915 1.16 ;
        RECT 1.915 1.04 2.155 1.195 ;
        RECT 0.65 1.075 0.8 1.435 ;
        RECT 0.435 1.075 0.8 1.195 ;
    END
  END B0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.42 1.175 4.57 1.435 ;
        RECT 4.195 1.175 4.57 1.315 ;
        RECT 4.195 1.075 4.315 1.315 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.595 1.045 3.835 1.195 ;
        RECT 3.495 0.94 3.755 1.12 ;
    END
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1072 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.075 1.555 3.195 2.21 ;
        RECT 0.07 1.555 3.195 1.675 ;
        RECT 2.395 0.735 2.635 0.855 ;
        RECT 0.195 0.785 2.515 0.905 ;
        RECT 2.235 1.555 2.355 2.21 ;
        RECT 1.395 1.555 1.515 2.21 ;
        RECT 0.915 0.735 1.155 0.905 ;
        RECT 0.555 1.555 0.675 2.21 ;
        RECT 0.195 0.785 0.315 1.675 ;
        RECT 0.07 1.465 0.22 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.495 -0.18 3.615 0.725 ;
        RECT 1.655 0.545 1.895 0.665 ;
        RECT 1.655 -0.18 1.775 0.665 ;
        RECT 0.275 0.545 0.515 0.665 ;
        RECT 0.275 -0.18 0.395 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 4.335 1.56 4.455 2.79 ;
        RECT 3.495 1.56 3.615 2.79 ;
        RECT 2.655 1.795 2.775 2.79 ;
        RECT 1.815 1.795 1.935 2.79 ;
        RECT 0.975 1.795 1.095 2.79 ;
        RECT 0.135 1.845 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.255 0.955 4.075 0.955 4.075 1.555 4.035 1.555 4.035 2.21 3.915 2.21 3.915 1.435 1.295 1.435 1.295 1.4 1.175 1.4 1.175 1.28 1.415 1.28 1.415 1.315 2.435 1.315 2.435 1.28 2.675 1.28 2.675 1.315 3.955 1.315 3.955 0.835 4.135 0.835 4.135 0.675 4.255 0.675 ;
  END
END OAI2BB1X4

MACRO OA22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 1.42 1.195 1.66 ;
        RECT 0.94 1.465 1.135 1.725 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.28 0.51 1.74 ;
        RECT 0.38 1.28 0.5 1.76 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.28 0.82 1.715 ;
        RECT 0.65 1.31 0.8 1.725 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.46 1.96 1.725 ;
        RECT 1.555 1.46 1.96 1.58 ;
        RECT 1.555 1.42 1.675 1.665 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.65 2.745 0.77 ;
        RECT 2.215 1.005 2.54 1.145 ;
        RECT 2.39 0.65 2.54 1.145 ;
        RECT 2.215 1.005 2.335 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.985 -0.18 3.105 0.64 ;
        RECT 2.085 -0.18 2.205 0.53 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.635 1.56 2.755 2.79 ;
        RECT 1.795 1.845 1.915 2.79 ;
        RECT 0.22 1.88 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.095 1.3 1.435 1.3 1.435 1.965 0.915 1.965 0.915 1.845 1.315 1.845 1.315 0.8 1.395 0.8 1.395 0.68 1.515 0.68 1.515 0.92 1.435 0.92 1.435 1.18 2.095 1.18 ;
      POLYGON 1.935 0.92 1.815 0.92 1.815 0.56 1.095 0.56 1.095 1.16 0.195 1.16 0.195 0.86 0.075 0.86 0.075 0.74 0.315 0.74 0.315 1.04 0.975 1.04 0.975 0.44 1.935 0.44 ;
  END
END OA22X2

MACRO NAND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X8 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.555 1.05 8.795 1.17 ;
        RECT 8.555 0.73 8.675 1.17 ;
        RECT 5.64 0.73 8.675 0.85 ;
        RECT 6.315 1.03 6.555 1.15 ;
        RECT 6.435 0.73 6.555 1.15 ;
        RECT 1.55 0.725 5.76 0.845 ;
        RECT 4.05 1.03 4.29 1.15 ;
        RECT 4.05 0.725 4.17 1.15 ;
        RECT 1.43 1.035 1.67 1.155 ;
        RECT 1.55 0.725 1.67 1.155 ;
        RECT 1.52 0.885 1.67 1.155 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.765 1.03 8.435 1.15 ;
        RECT 8.135 1.03 8.395 1.38 ;
        RECT 6.97 0.97 7.885 1.09 ;
        RECT 6.705 1.05 7.195 1.17 ;
        RECT 5.91 1.27 6.825 1.39 ;
        RECT 6.705 1.05 6.825 1.39 ;
        RECT 5.91 1.11 6.03 1.39 ;
        RECT 5.38 1.11 6.03 1.23 ;
        RECT 5.38 0.965 5.5 1.23 ;
        RECT 4.78 0.965 5.5 1.085 ;
        RECT 4.41 1.105 4.9 1.225 ;
        RECT 4.78 0.965 4.9 1.225 ;
        RECT 3.81 1.27 4.53 1.39 ;
        RECT 4.41 1.105 4.53 1.39 ;
        RECT 3.81 1.05 3.93 1.39 ;
        RECT 3.015 1.05 3.93 1.17 ;
        RECT 2.22 0.965 3.135 1.085 ;
        RECT 1.935 1.045 2.34 1.165 ;
        RECT 1.935 1.045 2.095 1.285 ;
        RECT 1.14 1.275 2.055 1.395 ;
        RECT 1.14 1.055 1.26 1.395 ;
        RECT 0.755 1.055 1.26 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.355 1.21 7.595 1.33 ;
        RECT 6.995 1.29 7.475 1.41 ;
        RECT 3.55 1.51 7.115 1.63 ;
        RECT 6.995 1.29 7.115 1.63 ;
        RECT 5.14 1.205 5.26 1.63 ;
        RECT 5.02 1.205 5.26 1.325 ;
        RECT 3.55 1.29 3.67 1.63 ;
        RECT 2.49 1.29 3.67 1.41 ;
        RECT 2.635 1.205 2.875 1.41 ;
        RECT 0.9 1.515 2.61 1.635 ;
        RECT 2.49 1.29 2.61 1.635 ;
        RECT 0.9 1.295 1.02 1.635 ;
        RECT 0.39 1.295 1.02 1.415 ;
        RECT 0.39 0.885 0.51 1.415 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.194 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.955 1.47 9.075 2.21 ;
        RECT 8.77 1.465 9.035 1.875 ;
        RECT 8.915 0.485 9.035 1.875 ;
        RECT 1.435 0.485 9.035 0.605 ;
        RECT 0.555 1.755 9.075 1.875 ;
        RECT 8.115 1.5 8.235 2.21 ;
        RECT 7.275 1.53 7.395 2.21 ;
        RECT 6.435 1.75 6.555 2.21 ;
        RECT 5.595 1.75 5.715 2.21 ;
        RECT 4.755 1.75 4.875 2.21 ;
        RECT 3.915 1.75 4.035 2.21 ;
        RECT 3.075 1.53 3.195 2.21 ;
        RECT 2.235 1.755 2.355 2.21 ;
        RECT 1.395 1.755 1.515 2.21 ;
        RECT 0.555 1.535 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 7.635 -0.18 7.875 0.365 ;
        RECT 5.25 -0.18 5.49 0.365 ;
        RECT 2.455 -0.18 2.695 0.365 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 8.475 1.995 8.715 2.15 ;
        RECT 8.475 1.995 8.595 2.79 ;
        RECT 7.635 1.995 7.875 2.15 ;
        RECT 7.635 1.995 7.755 2.79 ;
        RECT 6.795 1.995 7.035 2.15 ;
        RECT 6.795 1.995 6.915 2.79 ;
        RECT 5.955 1.995 6.195 2.15 ;
        RECT 5.955 1.995 6.075 2.79 ;
        RECT 5.115 1.995 5.355 2.15 ;
        RECT 5.115 1.995 5.235 2.79 ;
        RECT 4.275 1.995 4.515 2.15 ;
        RECT 4.275 1.995 4.395 2.79 ;
        RECT 3.435 1.995 3.675 2.15 ;
        RECT 3.435 1.995 3.555 2.79 ;
        RECT 2.595 1.995 2.835 2.15 ;
        RECT 2.595 1.995 2.715 2.79 ;
        RECT 1.755 1.995 1.995 2.15 ;
        RECT 1.755 1.995 1.875 2.79 ;
        RECT 0.915 1.995 1.155 2.15 ;
        RECT 0.915 1.995 1.035 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
END NAND3X8

MACRO SDFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX4 0 0 ;
  SIZE 13.63 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.615 0.36 1.735 1.53 ;
        RECT 0.895 0.36 1.735 0.48 ;
        RECT 0.92 0.92 1.235 1.04 ;
        RECT 0.39 0.9 1.04 1.02 ;
        RECT 0.895 0.36 1.015 1.02 ;
        RECT 0.36 1.175 0.51 1.435 ;
        RECT 0.39 0.9 0.51 1.435 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.16 0.835 1.53 ;
        RECT 0.65 1.14 0.8 1.53 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.29 2.25 1.435 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.935 1.29 2.055 1.53 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.06 2.54 1.53 ;
        RECT 2.37 0.96 2.49 1.46 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.835 1 8.955 1.24 ;
        RECT 7.795 1 8.955 1.12 ;
        RECT 7.915 0.57 8.035 1.12 ;
        RECT 7.195 0.57 8.035 0.69 ;
        RECT 7.195 0.38 7.315 0.69 ;
        RECT 6.295 0.38 7.315 0.5 ;
        RECT 5.385 1.24 6.415 1.36 ;
        RECT 6.295 0.38 6.415 1.36 ;
        RECT 6.245 0.94 6.415 1.36 ;
        RECT 6.105 0.94 6.415 1.09 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.715 1.44 10.835 2.21 ;
        RECT 10.535 1.44 10.835 1.56 ;
        RECT 9.475 0.68 10.675 0.8 ;
        RECT 9.93 1.32 10.655 1.44 ;
        RECT 9.93 1.175 10.08 1.44 ;
        RECT 9.93 0.68 10.05 1.56 ;
        RECT 9.875 1.44 9.995 2.21 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.395 0.68 12.595 0.8 ;
        RECT 12.395 1.44 12.515 2.21 ;
        RECT 12.215 1.44 12.515 1.56 ;
        RECT 11.67 1.32 12.335 1.44 ;
        RECT 11.67 1.175 11.82 1.44 ;
        RECT 11.67 0.68 11.79 1.56 ;
        RECT 11.555 1.44 11.675 2.21 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.63 0.18 ;
        RECT 12.835 -0.18 13.075 0.32 ;
        RECT 11.875 -0.18 12.115 0.32 ;
        RECT 10.915 -0.18 11.155 0.32 ;
        RECT 9.955 -0.18 10.195 0.32 ;
        RECT 8.995 -0.18 9.235 0.32 ;
        RECT 7.595 0.33 7.835 0.45 ;
        RECT 7.595 -0.18 7.715 0.45 ;
        RECT 5.875 0.68 6.175 0.8 ;
        RECT 6.055 -0.18 6.175 0.8 ;
        RECT 2.955 -0.18 3.075 0.92 ;
        RECT 1.895 -0.18 2.015 0.78 ;
        RECT 0.555 -0.18 0.675 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.63 2.79 ;
        RECT 12.815 1.56 12.935 2.79 ;
        RECT 11.975 1.56 12.095 2.79 ;
        RECT 11.135 1.56 11.255 2.79 ;
        RECT 10.295 1.56 10.415 2.79 ;
        RECT 9.455 1.56 9.575 2.79 ;
        RECT 8.315 1.72 8.435 2.79 ;
        RECT 7.415 1.72 7.655 2.09 ;
        RECT 7.415 1.72 7.535 2.79 ;
        RECT 5.935 2.17 6.055 2.79 ;
        RECT 5.815 2.17 6.055 2.29 ;
        RECT 4.735 2.2 4.975 2.79 ;
        RECT 3.14 2 3.26 2.79 ;
        RECT 2.095 1.89 2.215 2.79 ;
        RECT 0.635 1.89 0.755 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.495 0.86 13.355 0.86 13.355 2.21 13.235 2.21 13.235 1.44 12.655 1.44 12.655 1.2 12.775 1.2 12.775 1.32 13.235 1.32 13.235 0.74 13.375 0.74 13.375 0.62 13.495 0.62 ;
      POLYGON 13.095 1.2 12.975 1.2 12.975 0.56 10.915 0.56 10.915 1.06 10.895 1.06 10.895 1.18 10.775 1.18 10.775 0.94 10.795 0.94 10.795 0.56 8.475 0.56 8.475 0.76 8.355 0.76 8.355 0.44 13.095 0.44 ;
      POLYGON 9.335 1.6 8.855 1.6 8.855 2.15 8.735 2.15 8.735 1.6 8.015 1.6 8.015 2.15 7.895 2.15 7.895 1.6 7.315 1.6 7.315 1.31 7.435 1.31 7.435 1.48 9.215 1.48 9.215 1.22 9.335 1.22 ;
      POLYGON 8.375 1.36 7.555 1.36 7.555 0.93 6.915 0.93 6.915 1.81 6.955 1.81 6.955 1.93 6.715 1.93 6.715 1.81 6.795 1.81 6.795 0.74 6.955 0.74 6.955 0.62 7.075 0.62 7.075 0.81 7.675 0.81 7.675 1.24 8.375 1.24 ;
      POLYGON 7.275 1.17 7.195 1.17 7.195 2.17 6.815 2.17 6.815 2.25 6.575 2.25 6.575 2.17 6.175 2.17 6.175 2.05 5.695 2.05 5.695 2.2 5.095 2.2 5.095 2.08 4.345 2.08 4.345 2.06 4.335 2.06 4.335 2 3.42 2 3.42 1.88 4.345 1.88 4.345 1.82 4.465 1.82 4.465 1.96 5.215 1.96 5.215 2.08 5.575 2.08 5.575 1.93 6.295 1.93 6.295 2.05 7.075 2.05 7.075 1.17 7.035 1.17 7.035 1.05 7.275 1.05 ;
      POLYGON 6.655 1.69 6.535 1.69 6.535 1.81 6.295 1.81 6.295 1.6 5.085 1.6 5.085 1.31 5.205 1.31 5.205 1.48 6.535 1.48 6.535 0.62 6.655 0.62 ;
      POLYGON 5.985 1.12 4.845 1.12 4.845 1.22 4.485 1.22 4.485 1.58 4.305 1.58 4.305 1.7 4.185 1.7 4.185 1.46 4.365 1.46 4.365 1.1 4.725 1.1 4.725 0.62 4.845 0.62 4.845 1 5.985 1 ;
      POLYGON 5.935 0.48 4.415 0.48 4.415 0.5 4.15 0.5 4.15 0.74 3.885 0.74 3.885 0.98 4.005 0.98 4.005 1.1 3.765 1.1 3.765 0.98 3.555 0.98 3.555 1.52 3.315 1.52 3.315 1.4 3.435 1.4 3.435 0.86 3.315 0.86 3.315 0.74 3.555 0.74 3.555 0.86 3.765 0.86 3.765 0.62 4.03 0.62 4.03 0.38 4.295 0.38 4.295 0.36 5.935 0.36 ;
      POLYGON 5.455 1.96 5.335 1.96 5.335 1.84 4.605 1.84 4.605 1.34 4.725 1.34 4.725 1.72 5.455 1.72 ;
      POLYGON 4.425 0.98 4.245 0.98 4.245 1.34 3.885 1.34 3.885 1.76 3.02 1.76 3.02 2.25 2.335 2.25 2.335 1.77 1.8 1.77 1.8 1.89 1.535 1.89 1.535 2.01 1.415 2.01 1.415 1.89 1.375 1.89 1.375 0.72 1.135 0.72 1.135 0.6 1.495 0.6 1.495 1.77 1.68 1.77 1.68 1.65 2.455 1.65 2.455 2.13 2.9 2.13 2.9 1.64 3.765 1.64 3.765 1.22 4.125 1.22 4.125 0.86 4.305 0.86 4.305 0.62 4.425 0.62 ;
      POLYGON 3.275 1.2 2.78 1.2 2.78 1.77 2.695 1.77 2.695 2.01 2.575 2.01 2.575 1.65 2.66 1.65 2.66 0.84 2.315 0.84 2.315 0.54 2.435 0.54 2.435 0.72 2.78 0.72 2.78 1.08 3.275 1.08 ;
      POLYGON 1.255 1.77 0.335 1.77 0.335 2.01 0.215 2.01 0.215 1.89 0.12 1.89 0.12 0.935 0.135 0.935 0.135 0.54 0.255 0.54 0.255 1.055 0.24 1.055 0.24 1.65 1.135 1.65 1.135 1.45 1.255 1.45 ;
  END
END SDFFRX4

MACRO TLATSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX1 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.52 ;
        RECT 1.945 1.26 2.25 1.43 ;
    END
  END SN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.2 3.005 1.45 ;
        RECT 2.625 1.2 2.885 1.47 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.16 3.845 1.41 ;
        RECT 3.495 1.14 3.755 1.41 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 1.28 5.835 1.735 ;
        RECT 5.715 1.26 5.835 1.735 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2888 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 0.92 ;
        RECT 1.285 0.8 1.405 2.21 ;
        RECT 1.23 1.465 1.405 1.725 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 5.955 -0.18 6.075 0.78 ;
        RECT 4.025 0.42 4.265 0.54 ;
        RECT 4.145 -0.18 4.265 0.54 ;
        RECT 1.785 -0.18 1.905 0.73 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 5.875 2.2 6.115 2.79 ;
        RECT 4.305 2.01 4.425 2.79 ;
        RECT 3.465 2.23 3.585 2.79 ;
        RECT 2.605 2.23 2.725 2.79 ;
        RECT 1.705 1.59 1.825 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.535 1.84 6.415 1.84 6.415 1.72 6.375 1.72 6.375 1.02 5.595 1.02 5.595 1.14 5.475 1.14 5.475 0.9 6.375 0.9 6.375 0.54 6.495 0.54 6.495 1.6 6.535 1.6 ;
      POLYGON 6.475 2.22 6.235 2.22 6.235 2.08 5.555 2.08 5.555 2.22 5.315 2.22 5.315 2.08 4.995 2.08 4.995 1.04 4.875 1.04 4.875 1.02 3.375 1.02 3.375 1.71 3.105 1.71 3.105 1.83 2.985 1.83 2.985 1.59 3.255 1.59 3.255 0.6 3.565 0.6 3.565 0.72 3.375 0.72 3.375 0.9 5.115 0.9 5.115 1.96 6.355 1.96 6.355 2.1 6.475 2.1 ;
      POLYGON 5.355 1.84 5.235 1.84 5.235 0.78 3.73 0.78 3.73 0.48 2.79 0.48 2.79 0.54 2.285 0.54 2.285 0.42 2.67 0.42 2.67 0.36 3.85 0.36 3.85 0.66 5.215 0.66 5.215 0.54 5.335 0.54 5.335 0.66 5.355 0.66 ;
      POLYGON 4.875 1.8 4.755 1.8 4.755 1.89 3.765 1.89 3.765 1.77 4.635 1.77 4.635 1.68 4.875 1.68 ;
      POLYGON 4.225 1.65 3.645 1.65 3.645 2.07 2.125 2.07 2.125 1.64 2.37 1.64 2.37 1.055 1.725 1.055 1.725 1.26 1.605 1.26 1.605 0.935 2.485 0.935 2.485 0.68 2.605 0.68 2.605 1.055 2.49 1.055 2.49 1.76 2.245 1.76 2.245 1.95 3.525 1.95 3.525 1.53 4.105 1.53 4.105 1.27 4.225 1.27 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END TLATSRX1

MACRO OAI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X1 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.12 1.96 1.435 ;
        RECT 1.74 0.96 1.86 1.27 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 1.035 1.38 1.47 ;
        RECT 1.21 1.01 1.33 1.47 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.165 1.09 1.435 ;
        RECT 0.815 1.165 1.09 1.285 ;
        RECT 0.815 1.035 0.935 1.285 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3284 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.3 0.675 2.19 ;
        RECT 0.255 1.3 0.675 1.42 ;
        RECT 0.255 0.6 0.375 1.42 ;
        RECT 0.07 0.885 0.375 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 0.975 -0.18 1.095 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 2.23 1.895 2.79 ;
        RECT 0.975 1.59 1.095 2.79 ;
        RECT 0.135 1.54 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.81 0.84 1.62 0.84 1.62 1.71 1.515 1.71 1.515 1.83 1.395 1.83 1.395 1.59 1.5 1.59 1.5 0.89 0.615 0.89 0.615 1.18 0.495 1.18 0.495 0.77 1.5 0.77 1.5 0.72 1.69 0.72 1.69 0.6 1.81 0.6 ;
  END
END OAI2BB1X1

MACRO DLY4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X1 0 0 ;
  SIZE 10.15 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.64 1.165 9.79 1.615 ;
        RECT 9.64 1.165 9.76 1.64 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.875 0.94 1.145 1.09 ;
        RECT 0.875 0.68 0.995 1.99 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.15 0.18 ;
        RECT 9.475 -0.18 9.595 0.765 ;
        RECT 9.075 -0.18 9.195 1.005 ;
        RECT 8.975 0.885 9.095 1.48 ;
        RECT 7.605 -0.18 7.725 0.38 ;
        RECT 6.715 1.3 6.955 1.42 ;
        RECT 6.835 -0.18 6.955 1.42 ;
        RECT 5.875 1.24 6.115 1.36 ;
        RECT 5.965 -0.18 6.085 1.36 ;
        RECT 5.325 -0.18 5.445 0.38 ;
        RECT 4.585 -0.18 4.705 1.09 ;
        RECT 4.555 0.97 4.675 1.77 ;
        RECT 3.655 1.59 3.935 1.71 ;
        RECT 3.655 -0.18 3.775 1.71 ;
        RECT 3.195 -0.18 3.315 0.53 ;
        RECT 2.725 1.2 2.845 1.44 ;
        RECT 2.685 -0.18 2.805 1.32 ;
        RECT 1.885 -0.18 2.005 0.92 ;
        RECT 0.395 -0.18 0.515 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.15 2.79 ;
        RECT 9.475 1.76 9.595 2.79 ;
        RECT 8.205 1 8.325 1.24 ;
        RECT 7.075 1.04 8.325 1.16 ;
        RECT 7.695 2.2 7.815 2.79 ;
        RECT 7.295 1.04 7.415 2.79 ;
        RECT 5.315 2.2 5.555 2.79 ;
        RECT 4.295 1.04 4.415 2.79 ;
        RECT 4.175 1.04 4.415 1.16 ;
        RECT 3.135 2.08 3.375 2.2 ;
        RECT 3.235 2.08 3.355 2.79 ;
        RECT 2.325 1.04 2.565 1.18 ;
        RECT 1.505 1.04 2.565 1.16 ;
        RECT 1.505 2.28 1.925 2.79 ;
        RECT 1.505 1.04 1.625 2.79 ;
        RECT 0.455 1.34 0.575 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.03 1.88 10.015 1.88 10.015 2 9.895 2 9.895 1.76 9.91 1.76 9.91 1.045 9.315 1.045 9.315 0.925 9.895 0.925 9.895 0.525 10.015 0.525 10.015 0.805 10.03 0.805 ;
      POLYGON 8.955 0.765 8.855 0.765 8.855 1.64 8.955 1.64 8.955 1.88 8.835 1.88 8.835 1.76 8.735 1.76 8.735 0.645 8.835 0.645 8.835 0.525 8.8 0.525 8.8 0.52 7.885 0.52 7.885 0.4 8.92 0.4 8.92 0.405 8.955 0.405 ;
      POLYGON 8.565 1.48 8.485 1.48 8.485 1.8 8.365 1.8 8.365 1.48 7.535 1.48 7.535 1.3 7.775 1.3 7.775 1.36 8.445 1.36 8.445 0.66 8.565 0.66 ;
      POLYGON 7.175 1.84 5.295 1.84 5.295 1.75 5.275 1.75 5.275 1.51 5.295 1.51 5.295 0.5 5.605 0.5 5.605 0.4 5.845 0.4 5.845 0.62 5.415 0.62 5.415 1.72 6.475 1.72 6.475 0.78 6.595 0.78 6.595 0.66 6.715 0.66 6.715 0.9 6.595 0.9 6.595 1.72 7.175 1.72 ;
      POLYGON 6.355 1.6 5.535 1.6 5.535 1.48 6.235 1.48 6.235 1.12 6.205 1.12 6.205 0.66 6.325 0.66 6.325 1 6.355 1 ;
      POLYGON 6.255 2.08 5.035 2.08 5.035 1.09 4.945 1.09 4.945 0.48 4.825 0.48 4.825 0.36 5.065 0.36 5.065 0.97 5.155 0.97 5.155 1.96 6.255 1.96 ;
      POLYGON 4.915 2.01 4.795 2.01 4.795 2.13 4.675 2.13 4.675 1.89 4.795 1.89 4.795 1.21 4.915 1.21 ;
      POLYGON 4.465 0.84 4.225 0.84 4.225 0.48 4.145 0.48 4.145 0.36 4.385 0.36 4.385 0.48 4.345 0.48 4.345 0.72 4.465 0.72 ;
      POLYGON 4.175 1.97 4.015 1.97 4.015 2.09 3.895 2.09 3.895 1.97 3.735 1.97 3.735 1.96 2.795 1.96 2.795 2.16 2.025 2.16 2.025 2.04 2.675 2.04 2.675 1.84 3.855 1.84 3.855 1.85 4.055 1.85 4.055 1.47 3.935 1.47 3.935 0.86 3.895 0.86 3.895 0.62 4.015 0.62 4.015 0.74 4.055 0.74 4.055 1.35 4.175 1.35 ;
      POLYGON 3.085 1.72 2.525 1.72 2.525 1.68 2.445 1.68 2.445 1.42 1.745 1.42 1.745 1.28 1.985 1.28 1.985 1.3 2.565 1.3 2.565 1.56 2.965 1.56 2.965 0.92 2.925 0.92 2.925 0.68 3.045 0.68 3.045 0.8 3.085 0.8 ;
      POLYGON 1.585 0.92 1.385 0.92 1.385 1.78 1.265 1.78 1.265 0.8 1.465 0.8 1.465 0.68 1.43 0.68 1.43 0.56 0.755 0.56 0.755 1.18 0.515 1.18 0.515 1.06 0.635 1.06 0.635 0.44 1.55 0.44 1.55 0.56 1.585 0.56 ;
  END
END DLY4X1

MACRO ADDFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX4 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.035 0.82 7.495 0.94 ;
        RECT 5.175 0.82 5.415 1.09 ;
        RECT 4.055 0.78 5.155 0.9 ;
        RECT 4.075 0.65 4.335 0.9 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 0.94 8.395 1.25 ;
        RECT 8.135 0.94 8.395 1.16 ;
        RECT 7.655 1.04 8.395 1.16 ;
        RECT 5.535 1.06 7.775 1.18 ;
        RECT 4.795 1.21 5.655 1.33 ;
        RECT 5.535 1.06 5.655 1.33 ;
        RECT 4.795 1.02 4.915 1.33 ;
        RECT 3.735 1.02 4.915 1.14 ;
        RECT 2.675 0.98 3.855 1.1 ;
        RECT 2.675 0.98 2.795 1.24 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.895 1.28 8.135 1.4 ;
        RECT 5.775 1.3 8.015 1.42 ;
        RECT 4.42 1.45 5.895 1.57 ;
        RECT 5.775 1.3 5.895 1.57 ;
        RECT 4.42 1.28 4.675 1.57 ;
        RECT 4.42 1.28 4.57 1.725 ;
        RECT 4.05 1.28 4.675 1.4 ;
        RECT 3.135 1.26 4.17 1.34 ;
        RECT 3.255 1.28 4.675 1.38 ;
        RECT 3.135 1.22 3.375 1.34 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.32 1.555 2.21 ;
        RECT 1.435 0.67 1.555 0.96 ;
        RECT 0.555 1.32 1.555 1.44 ;
        RECT 0.555 0.84 1.555 0.96 ;
        RECT 0.595 1.32 0.715 2.21 ;
        RECT 0.595 0.67 0.715 0.96 ;
        RECT 0.555 0.79 0.675 1.44 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.735 0.885 10.08 1.145 ;
        RECT 8.855 1.32 9.855 1.44 ;
        RECT 9.735 0.76 9.855 1.44 ;
        RECT 9.695 1.32 9.815 2.21 ;
        RECT 8.855 0.76 9.855 0.88 ;
        RECT 9.695 0.59 9.815 0.88 ;
        RECT 8.855 1.32 8.975 2.21 ;
        RECT 8.855 0.59 8.975 0.88 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 10.115 -0.18 10.235 0.64 ;
        RECT 9.275 -0.18 9.395 0.64 ;
        RECT 8.375 0.46 8.615 0.58 ;
        RECT 8.375 -0.18 8.495 0.58 ;
        RECT 5.935 0.34 6.175 0.46 ;
        RECT 5.935 -0.18 6.055 0.46 ;
        RECT 5.095 -0.18 5.215 0.64 ;
        RECT 2.815 -0.18 3.055 0.38 ;
        RECT 1.855 -0.18 1.975 0.72 ;
        RECT 1.015 -0.18 1.135 0.72 ;
        RECT 0.175 -0.18 0.295 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 10.115 1.56 10.235 2.79 ;
        RECT 9.275 1.56 9.395 2.79 ;
        RECT 8.375 2.02 8.615 2.15 ;
        RECT 8.375 2.02 8.495 2.79 ;
        RECT 5.935 2.17 6.175 2.79 ;
        RECT 4.975 2.17 5.215 2.79 ;
        RECT 2.875 2.1 2.995 2.79 ;
        RECT 1.795 2.03 2.035 2.15 ;
        RECT 1.795 2.03 1.915 2.79 ;
        RECT 1.015 1.56 1.135 2.79 ;
        RECT 0.175 1.56 0.295 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.615 1.12 8.635 1.12 8.635 1.9 7.655 1.9 7.655 2.15 7.415 2.15 7.415 1.9 7.255 1.9 7.255 2.15 7.015 2.15 7.015 1.88 7.135 1.88 7.135 1.78 8.515 1.78 8.515 0.82 8.135 0.82 8.135 0.7 6.835 0.7 6.835 0.58 7.515 0.58 7.515 0.5 7.755 0.5 7.755 0.58 8.255 0.58 8.255 0.7 8.635 0.7 8.635 1 9.615 1 ;
      POLYGON 7.335 1.66 6.895 1.66 6.895 2.05 4.455 2.05 4.455 2.21 4.335 2.21 4.335 2.05 3.895 2.05 3.895 2.15 3.775 2.15 3.775 2.05 3.685 2.05 3.685 1.98 2.36 1.98 2.36 1.91 2.095 1.91 2.095 1.2 0.795 1.2 0.795 1.08 2.095 1.08 2.095 0.5 3.775 0.5 3.775 0.41 4.575 0.41 4.575 0.65 4.455 0.65 4.455 0.53 3.895 0.53 3.895 0.74 3.775 0.74 3.775 0.62 2.215 0.62 2.215 1.79 2.48 1.79 2.48 1.86 3.775 1.86 3.775 1.5 3.895 1.5 3.895 1.93 4.335 1.93 4.335 1.845 4.455 1.845 4.455 1.93 6.775 1.93 6.775 1.54 7.335 1.54 ;
      RECT 5.455 0.58 6.655 0.7 ;
      POLYGON 6.655 1.81 5.455 1.81 5.455 1.69 6.415 1.69 6.415 1.62 6.655 1.62 ;
      RECT 2.335 0.74 3.535 0.86 ;
      POLYGON 3.475 1.74 3.355 1.74 3.355 1.62 2.515 1.62 2.515 1.67 2.395 1.67 2.395 1.34 2.515 1.34 2.515 1.5 3.475 1.5 ;
  END
END ADDFX4

MACRO CLKAND2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X12 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.255 1 3.375 1.24 ;
        RECT 0.68 1 3.375 1.12 ;
        RECT 1.99 1 2.23 1.195 ;
        RECT 0.65 1.075 0.8 1.435 ;
        RECT 0.435 1.075 0.8 1.195 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.28 4.255 1.4 ;
        RECT 1.27 1.36 3.755 1.48 ;
        RECT 3.495 1.23 3.755 1.48 ;
        RECT 2.39 1.24 2.51 1.48 ;
        RECT 1.27 1.24 1.39 1.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.25 1.39 8.37 2.21 ;
        RECT 8.19 1.175 8.34 1.51 ;
        RECT 8.19 0.795 8.31 1.51 ;
        RECT 4.89 1.39 8.37 1.51 ;
        RECT 4.655 0.91 8.31 1.03 ;
        RECT 8.05 0.795 8.31 1.03 ;
        RECT 8.05 0.4 8.17 1.03 ;
        RECT 7.41 1.39 7.53 2.21 ;
        RECT 7.21 0.4 7.33 1.03 ;
        RECT 6.57 1.39 6.69 2.21 ;
        RECT 6.37 0.4 6.49 1.03 ;
        RECT 5.73 1.39 5.85 2.21 ;
        RECT 5.53 0.4 5.65 1.03 ;
        RECT 4.89 1.39 5.01 2.21 ;
        RECT 4.655 0.4 4.775 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.47 -0.18 8.59 0.915 ;
        RECT 7.63 -0.18 7.75 0.79 ;
        RECT 6.79 -0.18 6.91 0.79 ;
        RECT 5.95 -0.18 6.07 0.79 ;
        RECT 5.075 -0.18 5.195 0.79 ;
        RECT 4.235 -0.18 4.355 0.64 ;
        RECT 2.53 -0.18 2.65 0.64 ;
        RECT 0.99 -0.18 1.11 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.67 1.43 8.79 2.79 ;
        RECT 7.83 1.63 7.95 2.79 ;
        RECT 6.99 1.63 7.11 2.79 ;
        RECT 6.15 1.63 6.27 2.79 ;
        RECT 5.31 1.63 5.43 2.79 ;
        RECT 4.41 2.23 4.53 2.79 ;
        RECT 3.57 2.23 3.69 2.79 ;
        RECT 2.73 2.23 2.85 2.79 ;
        RECT 1.89 2.23 2.01 2.79 ;
        RECT 1.035 2.23 1.155 2.79 ;
        RECT 0.135 1.71 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.07 1.27 4.495 1.27 4.495 1.74 0.495 1.74 0.495 1.62 4.375 1.62 4.375 0.88 3.715 0.88 3.715 0.92 3.595 0.92 3.595 0.88 0.455 0.88 0.455 0.915 0.335 0.915 0.335 0.4 0.455 0.4 0.455 0.76 1.79 0.76 1.79 0.4 1.91 0.4 1.91 0.76 3.595 0.76 3.595 0.4 3.715 0.4 3.715 0.76 4.495 0.76 4.495 1.15 8.07 1.15 ;
  END
END CLKAND2X12

MACRO MXI3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3XL 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 1.465 1.575 1.585 ;
        RECT 0.305 1.52 1.455 1.62 ;
        RECT 0.355 1.5 1.575 1.585 ;
        RECT 0.305 1.52 0.565 1.67 ;
        RECT 0.355 1.38 0.475 1.67 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.23 1.115 1.35 ;
        RECT 0.595 1.23 0.855 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 1.395 2.54 1.725 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.515 1.42 4.475 1.54 ;
        RECT 3.515 1.23 3.755 1.54 ;
        RECT 3.515 1.18 3.635 1.54 ;
        RECT 3.495 1.23 3.755 1.38 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.965 1.175 5.175 1.435 ;
        RECT 4.965 1.04 5.15 1.435 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.665 0.68 5.785 1.6 ;
        RECT 5.58 0.885 5.785 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.245 -0.18 5.365 0.92 ;
        RECT 3.955 0.7 4.195 0.82 ;
        RECT 3.955 -0.18 4.075 0.82 ;
        RECT 2.255 0.7 2.495 0.82 ;
        RECT 2.255 -0.18 2.375 0.82 ;
        RECT 0.755 -0.18 0.875 0.87 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.125 2.1 5.365 2.22 ;
        RECT 5.125 2.1 5.245 2.79 ;
        RECT 3.695 2.265 3.935 2.79 ;
        RECT 2.315 1.845 2.435 2.79 ;
        RECT 0.875 1.845 0.995 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.705 1.98 5.005 1.98 5.005 2.145 3.83 2.145 3.83 2.1 3.035 2.1 3.035 1.86 2.855 1.86 2.855 0.7 3.135 0.7 3.135 0.82 2.975 0.82 2.975 1.74 3.155 1.74 3.155 1.98 3.95 1.98 3.95 2.025 4.885 2.025 4.885 1.86 5.705 1.86 ;
      POLYGON 4.945 0.92 4.845 0.92 4.845 1.3 4.825 1.3 4.825 1.6 4.705 1.6 4.705 1.3 3.875 1.3 3.875 1.18 4.725 1.18 4.725 0.8 4.825 0.8 4.825 0.68 4.945 0.68 ;
      POLYGON 4.555 1.06 3.375 1.06 3.375 1.5 3.395 1.5 3.395 1.665 4.295 1.665 4.295 1.785 4.415 1.785 4.415 1.905 4.175 1.905 4.175 1.785 3.275 1.785 3.275 1.62 3.215 1.62 3.215 1.585 3.095 1.585 3.095 1.465 3.255 1.465 3.255 0.58 2.855 0.58 2.855 0.48 2.735 0.48 2.735 0.36 2.975 0.36 2.975 0.46 3.505 0.46 3.505 0.94 4.435 0.94 4.435 0.64 4.555 0.64 ;
      POLYGON 2.595 1.275 2.475 1.275 2.475 1.265 2.195 1.265 2.195 1.865 1.855 1.865 1.855 1.905 1.615 1.905 1.615 1.785 1.735 1.785 1.735 1.745 2.075 1.745 2.075 1.265 2.015 1.265 2.015 0.82 1.395 0.82 1.395 0.7 2.135 0.7 2.135 1.145 2.475 1.145 2.475 1.035 2.595 1.035 ;
      POLYGON 1.955 1.625 1.835 1.625 1.835 1.505 1.695 1.505 1.695 1.16 1.235 1.16 1.235 1.11 0.185 1.11 0.185 1.79 0.575 1.79 0.575 2.03 0.455 2.03 0.455 1.91 0.065 1.91 0.065 0.87 0.275 0.87 0.275 0.64 0.395 0.64 0.395 0.99 1.815 0.99 1.815 1.385 1.955 1.385 ;
  END
END MXI3XL

MACRO NAND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X6 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.995 1.055 6.275 1.175 ;
        RECT 5.995 0.82 6.115 1.175 ;
        RECT 4.14 0.82 6.115 0.94 ;
        RECT 3.995 0.84 4.26 0.96 ;
        RECT 3.345 1.035 4.115 1.155 ;
        RECT 3.995 0.84 4.115 1.155 ;
        RECT 3.575 1.035 3.815 1.175 ;
        RECT 3.345 0.82 3.465 1.155 ;
        RECT 2.02 0.82 3.465 0.94 ;
        RECT 1.755 0.94 2.14 1.09 ;
        RECT 1.575 1.055 1.875 1.175 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.395 1.08 7.195 1.2 ;
        RECT 6.74 0.885 6.89 1.2 ;
        RECT 5.755 1.295 6.515 1.415 ;
        RECT 6.395 1.08 6.515 1.415 ;
        RECT 5.755 1.08 5.875 1.415 ;
        RECT 5.3 1.08 5.875 1.2 ;
        RECT 4.7 1.06 5.42 1.18 ;
        RECT 4.235 1.08 4.82 1.2 ;
        RECT 4.235 1.08 4.355 1.395 ;
        RECT 3.335 1.295 4.25 1.415 ;
        RECT 4.13 1.275 4.355 1.395 ;
        RECT 3.07 1.275 3.455 1.395 ;
        RECT 3.07 1.06 3.19 1.395 ;
        RECT 2.275 1.06 3.19 1.18 ;
        RECT 2.275 1.06 2.395 1.33 ;
        RECT 2.01 1.21 2.395 1.33 ;
        RECT 1.14 1.295 2.13 1.415 ;
        RECT 0.755 1.28 1.26 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.37 1.105 7.555 1.345 ;
        RECT 6.86 1.32 7.49 1.44 ;
        RECT 5.27 1.535 6.98 1.655 ;
        RECT 6.86 1.32 6.98 1.655 ;
        RECT 5.27 1.32 5.39 1.655 ;
        RECT 4.475 1.32 5.39 1.44 ;
        RECT 4.94 1.3 5.18 1.44 ;
        RECT 0.71 1.535 4.595 1.655 ;
        RECT 4.475 1.32 4.595 1.655 ;
        RECT 2.71 1.3 2.95 1.655 ;
        RECT 0.445 1.52 0.83 1.64 ;
        RECT 0.445 1.23 0.565 1.64 ;
        RECT 0.325 1.23 0.565 1.4 ;
        RECT 0.305 1.23 0.565 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.3781 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.775 7.795 1.895 ;
        RECT 7.675 0.58 7.795 1.895 ;
        RECT 7.61 1.465 7.795 1.895 ;
        RECT 1.295 0.58 7.795 0.7 ;
        RECT 7.275 1.56 7.395 2.21 ;
        RECT 6.435 1.775 6.555 2.21 ;
        RECT 6.235 0.4 6.355 0.915 ;
        RECT 5.595 1.775 5.715 2.21 ;
        RECT 4.755 1.56 4.875 2.21 ;
        RECT 3.915 1.775 4.035 2.21 ;
        RECT 3.755 0.4 3.875 0.915 ;
        RECT 3.075 1.775 3.195 2.21 ;
        RECT 2.235 1.775 2.355 2.21 ;
        RECT 1.395 1.775 1.515 2.21 ;
        RECT 1.295 0.4 1.415 0.92 ;
        RECT 0.555 1.775 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 5.075 0.34 5.315 0.46 ;
        RECT 5.075 -0.18 5.195 0.46 ;
        RECT 2.55 0.34 2.79 0.46 ;
        RECT 2.55 -0.18 2.67 0.46 ;
        RECT 0.335 -0.18 0.455 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.635 2.015 7.875 2.15 ;
        RECT 7.635 2.015 7.755 2.79 ;
        RECT 6.795 2.015 7.035 2.15 ;
        RECT 6.795 2.015 6.915 2.79 ;
        RECT 5.955 2.015 6.195 2.15 ;
        RECT 5.955 2.015 6.075 2.79 ;
        RECT 5.115 2.015 5.355 2.15 ;
        RECT 5.115 2.015 5.235 2.79 ;
        RECT 4.275 2.015 4.515 2.15 ;
        RECT 4.275 2.015 4.395 2.79 ;
        RECT 3.435 2.015 3.675 2.15 ;
        RECT 3.435 2.015 3.555 2.79 ;
        RECT 2.595 2.015 2.835 2.15 ;
        RECT 2.595 2.015 2.715 2.79 ;
        RECT 1.755 2.015 1.995 2.15 ;
        RECT 1.755 2.015 1.875 2.79 ;
        RECT 0.915 2.015 1.155 2.15 ;
        RECT 0.915 2.015 1.035 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND3X6

MACRO SDFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX2 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.87 2.885 1.1 ;
        RECT 2.695 0.87 2.815 1.28 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.76 2.05 6.325 2.17 ;
        RECT 4.76 1.87 4.88 2.17 ;
        RECT 4.685 1.435 4.805 1.99 ;
        RECT 4.13 1.435 4.805 1.555 ;
        RECT 4.13 1.175 4.28 1.555 ;
        RECT 3.945 1.17 4.25 1.29 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.77 1.175 9.085 1.32 ;
        RECT 8.965 1.08 9.085 1.32 ;
        RECT 8.77 1.175 8.92 1.435 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.025 1.3 10.305 1.42 ;
        RECT 9.875 1.81 10.145 1.96 ;
        RECT 10.025 1.3 10.145 1.96 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 1.175 10.66 1.435 ;
        RECT 9.785 1.06 10.63 1.18 ;
        RECT 10.51 1.055 10.63 1.435 ;
        RECT 9.785 1.06 9.905 1.5 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 0.885 1.38 1.145 ;
        RECT 1.035 1.4 1.315 1.52 ;
        RECT 1.195 0.59 1.315 1.52 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.885 2.25 1.145 ;
        RECT 1.995 1.4 2.235 1.52 ;
        RECT 2.035 0.59 2.155 1.52 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.225 -0.18 10.465 0.38 ;
        RECT 8.825 -0.18 8.945 0.92 ;
        RECT 5.925 -0.18 6.165 0.32 ;
        RECT 4.065 0.45 4.305 0.57 ;
        RECT 4.185 -0.18 4.305 0.57 ;
        RECT 2.455 -0.18 2.575 0.64 ;
        RECT 1.615 -0.18 1.735 0.64 ;
        RECT 0.775 -0.18 0.895 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.285 2.22 10.405 2.79 ;
        RECT 8.885 2.22 9.005 2.79 ;
        RECT 6.725 2.05 6.965 2.17 ;
        RECT 6.725 2.05 6.845 2.79 ;
        RECT 5.765 2.29 6.005 2.79 ;
        RECT 4.125 2.23 4.245 2.79 ;
        RECT 3.245 1.88 3.365 2.79 ;
        RECT 2.535 1.98 2.655 2.79 ;
        RECT 1.515 1.88 1.755 2 ;
        RECT 1.515 1.88 1.635 2.79 ;
        RECT 0.555 1.88 0.795 2 ;
        RECT 0.555 1.88 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.9 1.7 10.885 1.7 10.885 1.82 10.765 1.82 10.765 1.58 10.78 1.58 10.78 0.92 10.765 0.92 10.765 0.68 10.315 0.68 10.315 0.62 9.405 0.62 9.405 1.24 9.425 1.24 9.425 1.48 9.285 1.48 9.285 0.5 9.665 0.5 9.665 0.42 9.905 0.42 9.905 0.5 10.435 0.5 10.435 0.56 10.885 0.56 10.885 0.8 10.9 0.8 ;
      POLYGON 9.765 0.86 9.665 0.86 9.665 1.76 9.625 1.76 9.625 2 8.105 2 8.105 1.7 8.015 1.7 8.015 1.34 7.715 1.34 7.715 0.86 7.425 0.86 7.425 0.62 7.545 0.62 7.545 0.74 7.835 0.74 7.835 1.22 8.135 1.22 8.135 1.58 8.225 1.58 8.225 1.88 9.505 1.88 9.505 1.64 9.545 1.64 9.545 0.86 9.525 0.86 9.525 0.74 9.765 0.74 ;
      POLYGON 8.745 2.24 7.865 2.24 7.865 1.94 7.455 1.94 7.455 2.04 7.335 2.04 7.335 1.94 7.285 1.94 7.285 1.93 5.165 1.93 5.165 1.075 5.125 1.075 5.125 0.56 4.58 0.56 4.58 0.81 3.665 0.81 3.665 0.5 3.055 0.5 3.055 0.63 3.125 0.63 3.125 1.52 2.875 1.52 2.875 1.4 3.005 1.4 3.005 0.75 2.935 0.75 2.935 0.38 3.785 0.38 3.785 0.69 4.46 0.69 4.46 0.44 4.625 0.44 4.625 0.36 4.865 0.36 4.865 0.44 5.245 0.44 5.245 0.955 5.285 0.955 5.285 1.81 7.335 1.81 7.335 1.8 7.455 1.8 7.455 1.82 7.985 1.82 7.985 2.12 8.745 2.12 ;
      POLYGON 8.585 1.76 8.345 1.76 8.345 1.64 8.405 1.64 8.405 0.98 8.075 0.98 8.075 1.1 7.955 1.1 7.955 0.5 6.405 0.5 6.405 0.56 5.485 0.56 5.485 0.48 5.365 0.48 5.365 0.36 5.605 0.36 5.605 0.44 6.285 0.44 6.285 0.38 6.805 0.38 6.805 0.36 7.045 0.36 7.045 0.38 8.075 0.38 8.075 0.86 8.405 0.86 8.405 0.68 8.525 0.68 8.525 1.64 8.585 1.64 ;
      POLYGON 7.715 1.7 7.595 1.7 7.595 1.58 7.475 1.58 7.475 1.38 5.845 1.38 5.845 1.37 5.725 1.37 5.725 1.25 5.965 1.25 5.965 1.26 7.005 1.26 7.005 0.62 7.125 0.62 7.125 1.26 7.595 1.26 7.595 1.46 7.715 1.46 ;
      POLYGON 7.355 1.64 6.485 1.64 6.485 1.69 6.245 1.69 6.245 1.57 6.365 1.57 6.365 1.52 7.355 1.52 ;
      POLYGON 6.705 1.14 6.465 1.14 6.465 1.13 5.605 1.13 5.605 1.57 5.645 1.57 5.645 1.69 5.405 1.69 5.405 1.57 5.485 1.57 5.485 0.8 5.365 0.8 5.365 0.68 5.605 0.68 5.605 1.01 6.585 1.01 6.585 1.02 6.705 1.02 ;
      POLYGON 5.045 1.75 4.925 1.75 4.925 1.315 4.765 1.315 4.765 1.05 3.825 1.05 3.825 1.14 3.525 1.14 3.525 1.02 3.705 1.02 3.705 0.93 4.765 0.93 4.765 0.68 5.005 0.68 5.005 0.8 4.885 0.8 4.885 1.195 5.045 1.195 ;
      POLYGON 4.565 2.21 4.445 2.21 4.445 2.07 3.725 2.07 3.725 1.53 3.405 1.53 3.405 1.76 0.555 1.76 0.555 1 0.675 1 0.675 1.64 1.755 1.64 1.755 1.02 1.875 1.02 1.875 1.64 2.37 1.64 2.37 1 2.49 1 2.49 1.64 3.285 1.64 3.285 0.78 3.425 0.78 3.425 0.62 3.545 0.62 3.545 0.9 3.405 0.9 3.405 1.41 3.845 1.41 3.845 1.95 4.565 1.95 ;
      POLYGON 1.055 1.17 0.935 1.17 0.935 0.88 0.415 0.88 0.415 1.46 0.255 1.46 0.255 1.58 0.135 1.58 0.135 1.34 0.295 1.34 0.295 0.59 0.415 0.59 0.415 0.76 1.055 0.76 ;
  END
END SDFFRX2

MACRO MX3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X1 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.19 1.09 1.45 ;
        RECT 0.94 1.175 1.09 1.45 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.885 2.25 1.355 ;
        RECT 2.13 0.855 2.25 1.355 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.695 1.04 2.815 1.28 ;
        RECT 2.42 1.04 2.815 1.16 ;
        RECT 2.39 0.885 2.54 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.82 1.11 4.06 1.3 ;
        RECT 3.84 1.08 3.99 1.455 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.22 1.52 4.625 1.67 ;
        RECT 4.22 1.5 4.46 1.67 ;
        RECT 3.54 1.575 4.34 1.695 ;
        RECT 3.54 1.46 3.66 1.7 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 1.3 0.32 2.21 ;
        RECT 0.2 0.68 0.32 0.94 ;
        RECT 0.16 0.82 0.28 1.42 ;
        RECT 0.07 0.885 0.28 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.195 0.52 4.435 0.64 ;
        RECT 4.195 -0.18 4.315 0.64 ;
        RECT 2.975 -0.18 3.095 0.7 ;
        RECT 0.56 0.55 0.8 0.67 ;
        RECT 0.56 -0.18 0.68 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 4.04 1.9 4.16 2.79 ;
        RECT 2.76 1.9 2.88 2.79 ;
        RECT 0.62 1.72 0.74 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.865 1.91 4.58 1.91 4.58 2.03 4.46 2.03 4.46 1.79 4.745 1.79 4.745 0.96 3.7 0.96 3.7 1.34 3.295 1.34 3.295 1.48 3.175 1.48 3.175 1.22 3.58 1.22 3.58 0.84 4.745 0.84 4.745 0.7 4.675 0.7 4.675 0.46 4.795 0.46 4.795 0.58 4.865 0.58 ;
      POLYGON 3.795 0.64 3.46 0.64 3.46 1.1 3.055 1.1 3.055 1.66 3.42 1.66 3.42 1.82 3.52 1.82 3.52 2.06 3.4 2.06 3.4 1.94 3.3 1.94 3.3 1.78 2.13 1.78 2.13 1.9 1.86 1.9 1.86 0.6 2.1 0.6 2.1 0.72 1.98 0.72 1.98 1.66 2.935 1.66 2.935 0.98 3.34 0.98 3.34 0.52 3.795 0.52 ;
      POLYGON 2.675 0.7 2.555 0.7 2.555 0.48 1.74 0.48 1.74 2.02 2.34 2.02 2.34 1.9 2.46 1.9 2.46 2.14 1.62 2.14 1.62 1.64 1.45 1.64 1.45 1.4 1.62 1.4 1.62 1.04 1.5 1.04 1.5 0.92 1.62 0.92 1.62 0.36 2.675 0.36 ;
      POLYGON 1.5 0.72 1.38 0.72 1.38 1.055 1.33 1.055 1.33 1.78 1.5 1.78 1.5 1.9 1.21 1.9 1.21 1.055 0.7 1.055 0.7 1.18 0.4 1.18 0.4 1.06 0.58 1.06 0.58 0.935 1.26 0.935 1.26 0.6 1.5 0.6 ;
  END
END MX3X1

MACRO SDFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX1 0 0 ;
  SIZE 12.47 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.14 1.96 1.435 ;
        RECT 1.705 1.11 1.825 1.395 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.73 2.13 6.59 2.25 ;
        RECT 5.73 1.96 5.85 2.25 ;
        RECT 5.63 1.7 5.75 2.08 ;
        RECT 5.03 1.7 5.75 1.82 ;
        RECT 4.07 2.13 5.15 2.25 ;
        RECT 5.03 1.7 5.15 2.25 ;
        RECT 3.83 2.08 4.19 2.2 ;
        RECT 3.83 1.4 3.95 2.2 ;
        RECT 2.42 1.4 3.95 1.52 ;
        RECT 2.22 1.175 2.54 1.435 ;
        RECT 2.22 1.14 2.34 1.435 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 0.955 9.7 1.12 ;
        RECT 9.295 0.94 9.555 1.145 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.82 0.83 10.17 1.12 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.26 1.23 11.585 1.38 ;
        RECT 11.26 1.215 11.53 1.535 ;
        RECT 11.32 1.21 11.53 1.535 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.65 0.99 11.89 1.11 ;
        RECT 10.53 0.97 11.875 1.09 ;
        RECT 11.615 0.94 11.875 1.09 ;
        RECT 10.53 0.97 10.65 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 1.295 0.31 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.47 0.18 ;
        RECT 11.59 -0.18 11.71 0.82 ;
        RECT 10.07 -0.18 10.31 0.32 ;
        RECT 8.835 -0.18 9.075 0.32 ;
        RECT 7.01 0.49 7.25 0.61 ;
        RECT 7.01 -0.18 7.13 0.61 ;
        RECT 1.76 -0.18 2 0.32 ;
        RECT 0.555 -0.18 0.675 0.82 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.47 2.79 ;
        RECT 11.37 1.895 11.49 2.79 ;
        RECT 10.05 1.85 10.17 2.79 ;
        RECT 9.32 1.505 9.44 2.79 ;
        RECT 6.71 2.01 6.95 2.13 ;
        RECT 6.71 2.01 6.83 2.79 ;
        RECT 5.39 1.94 5.51 2.79 ;
        RECT 5.27 1.94 5.51 2.06 ;
        RECT 3.14 1.88 3.38 2 ;
        RECT 3.16 1.88 3.28 2.79 ;
        RECT 1.88 1.795 2 2.79 ;
        RECT 1.76 1.795 2 1.915 ;
        RECT 0.61 1.69 0.73 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.19 0.76 12.13 0.76 12.13 1.895 11.91 1.895 11.91 2.09 11.79 2.09 11.79 1.775 10.93 1.775 10.93 1.42 10.81 1.42 10.81 1.3 11.05 1.3 11.05 1.655 12.01 1.655 12.01 0.76 11.95 0.76 11.95 0.64 12.19 0.64 ;
      POLYGON 11.01 0.61 10.77 0.61 10.77 0.56 10.41 0.56 10.41 1.56 10.81 1.56 10.81 2.21 10.69 2.21 10.69 1.68 10.29 1.68 10.29 0.56 8.25 0.56 8.25 1.04 8.61 1.04 8.61 1.62 8.63 1.62 8.63 1.77 8.39 1.77 8.39 1.62 8.49 1.62 8.49 1.16 8.13 1.16 8.13 0.44 10.89 0.44 10.89 0.49 11.01 0.49 ;
      POLYGON 9.81 2.075 9.57 2.075 9.57 1.385 9.2 1.385 9.2 2.25 7.295 2.25 7.295 1.89 5.97 1.89 5.97 1.84 5.87 1.84 5.87 1.58 4.91 1.58 4.91 2.01 4.31 2.01 4.31 0.98 4.43 0.98 4.43 0.48 3.95 0.48 3.95 1.04 3.69 1.04 3.69 0.92 3.83 0.92 3.83 0.36 4.55 0.36 4.55 1.1 4.43 1.1 4.43 1.89 4.79 1.89 4.79 1.46 5.99 1.46 5.99 1.72 6.09 1.72 6.09 1.77 7.415 1.77 7.415 2.13 9.08 2.13 9.08 1.385 9.055 1.385 9.055 1.22 8.99 1.22 8.99 0.68 9.465 0.68 9.465 0.8 9.175 0.8 9.175 1.265 9.69 1.265 9.69 1.955 9.81 1.955 ;
      POLYGON 8.96 2.01 7.55 2.01 7.55 1.09 7.07 1.09 7.07 1.21 7 1.21 7 1.36 6.35 1.36 6.35 1.1 4.91 1.1 4.91 0.98 6.47 0.98 6.47 1.24 6.88 1.24 6.88 1.09 6.95 1.09 6.95 0.97 7.77 0.97 7.77 1.09 7.67 1.09 7.67 1.89 8.15 1.89 8.15 1.4 8.13 1.4 8.13 1.28 8.37 1.28 8.37 1.4 8.27 1.4 8.27 1.89 8.84 1.89 8.84 1.625 8.75 1.625 8.75 0.84 8.46 0.84 8.46 0.72 8.87 0.72 8.87 1.505 8.96 1.505 ;
      POLYGON 8.03 1.77 7.79 1.77 7.79 1.62 7.89 1.62 7.89 0.77 7.565 0.77 7.565 0.85 6.83 0.85 6.83 0.97 6.71 0.97 6.71 1.12 6.59 1.12 6.59 0.85 6.71 0.85 6.71 0.73 7.445 0.73 7.445 0.65 7.71 0.65 7.71 0.53 7.83 0.53 7.83 0.65 8.01 0.65 8.01 1.62 8.03 1.62 ;
      POLYGON 7.43 1.33 7.31 1.33 7.31 1.6 6.45 1.6 6.45 1.65 6.21 1.65 6.21 1.6 6.11 1.6 6.11 1.34 4.67 1.34 4.67 1.77 4.55 1.77 4.55 1.22 4.67 1.22 4.67 0.54 4.79 0.54 4.79 0.74 5.99 0.74 5.99 0.6 6.23 0.6 6.23 0.72 6.11 0.72 6.11 0.86 4.79 0.86 4.79 1.22 6.23 1.22 6.23 1.48 7.19 1.48 7.19 1.21 7.43 1.21 ;
      POLYGON 6.59 0.68 6.47 0.68 6.47 0.48 5.87 0.48 5.87 0.62 5.57 0.62 5.57 0.5 5.75 0.5 5.75 0.36 6.59 0.36 ;
      POLYGON 4.31 0.72 4.19 0.72 4.19 1.96 4.07 1.96 4.07 1.28 2.66 1.28 2.66 1.02 2.06 1.02 2.06 0.6 1.325 0.6 1.325 0.56 0.915 0.56 0.915 1.26 0.795 1.26 0.795 0.44 1.445 0.44 1.445 0.48 2.18 0.48 2.18 0.9 2.78 0.9 2.78 1.16 4.07 1.16 4.07 0.6 4.31 0.6 ;
      POLYGON 3.71 0.72 3.57 0.72 3.57 1.02 2.9 1.02 2.9 0.78 2.66 0.78 2.66 0.66 3.02 0.66 3.02 0.9 3.45 0.9 3.45 0.6 3.71 0.6 ;
      POLYGON 3.71 1.96 3.59 1.96 3.59 1.76 2.48 1.76 2.48 1.98 2.36 1.98 2.36 1.64 3.71 1.64 ;
      POLYGON 3.26 0.78 3.14 0.78 3.14 0.54 2.42 0.54 2.42 0.78 2.3 0.78 2.3 0.42 3.26 0.42 ;
      POLYGON 3.04 2.25 2.8 2.25 2.8 2.22 2.12 2.22 2.12 1.675 1.34 1.675 1.34 0.72 1.605 0.72 1.605 0.84 1.46 0.84 1.46 1.555 2.24 1.555 2.24 2.1 2.92 2.1 2.92 2.13 3.04 2.13 ;
      POLYGON 1.76 2.25 1.03 2.25 1.03 1.82 1.035 1.82 1.035 1.5 0.455 1.5 0.455 1.24 0.575 1.24 0.575 1.38 1.035 1.38 1.035 0.68 1.155 0.68 1.155 1.94 1.15 1.94 1.15 2.13 1.76 2.13 ;
  END
END SDFFSRHQX1

MACRO OAI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33XL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.37 1.14 2.61 1.345 ;
        RECT 2.39 1.08 2.54 1.475 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.105 2.25 1.56 ;
        RECT 2.1 1.08 2.22 1.56 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.175 1.38 1.675 ;
        RECT 1.23 1.175 1.38 1.645 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 1.24 0.54 1.62 ;
        RECT 0.07 1.315 0.54 1.435 ;
        RECT 0.07 1.06 0.22 1.435 ;
    END
  END A0
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.335 1.86 1.485 ;
        RECT 1.52 1.14 1.67 1.455 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.14 1.09 1.61 ;
        RECT 0.94 1.14 1.06 1.64 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2592 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.78 0.54 2.9 0.78 ;
        RECT 1.52 1.68 2.85 1.8 ;
        RECT 2.68 1.465 2.85 1.8 ;
        RECT 2.73 0.66 2.85 1.8 ;
        RECT 2 0.84 2.85 0.96 ;
        RECT 2 0.6 2.12 0.96 ;
        RECT 1.88 0.6 2.12 0.72 ;
        RECT 1.52 1.68 1.64 2.04 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 1.1 -0.18 1.22 0.78 ;
        RECT 0.26 -0.18 0.38 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.58 1.92 2.7 2.79 ;
        RECT 0.46 1.92 0.58 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.54 0.72 2.3 0.72 2.3 0.48 1.64 0.48 1.64 1.02 0.68 1.02 0.68 0.54 0.8 0.54 0.8 0.9 1.52 0.9 1.52 0.36 2.42 0.36 2.42 0.6 2.54 0.6 ;
  END
END OAI33XL

MACRO TLATSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX4 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7084 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.49 2.575 1.61 ;
        RECT 2.335 1.315 2.535 1.61 ;
        RECT 2.415 0.62 2.535 1.61 ;
        RECT 1.495 1.315 2.535 1.435 ;
        RECT 1.455 1.175 1.67 1.315 ;
        RECT 1.375 1.49 1.615 1.61 ;
        RECT 1.495 1.175 1.615 1.61 ;
        RECT 1.455 0.62 1.575 1.315 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.8 1.075 10.95 1.435 ;
        RECT 10.765 1.03 10.885 1.39 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.155 0.565 1.38 ;
        RECT 0.325 1.1 0.565 1.38 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.775 0.36 9.015 0.48 ;
        RECT 8.175 0.69 8.895 0.81 ;
        RECT 8.775 0.36 8.895 0.81 ;
        RECT 8.175 0.38 8.295 0.81 ;
        RECT 7.215 0.38 8.295 0.5 ;
        RECT 6.615 0.69 7.335 0.81 ;
        RECT 7.215 0.38 7.335 0.81 ;
        RECT 6.615 0.38 6.735 0.81 ;
        RECT 6.135 0.38 6.735 0.5 ;
        RECT 5.535 0.69 6.255 0.81 ;
        RECT 6.135 0.38 6.255 0.81 ;
        RECT 5.535 0.38 5.655 0.81 ;
        RECT 5.055 0.38 5.655 0.5 ;
        RECT 4.575 0.79 5.175 0.91 ;
        RECT 5.055 0.38 5.175 0.91 ;
        RECT 4.575 0.38 4.695 0.91 ;
        RECT 4.095 0.38 4.695 0.5 ;
        RECT 3.615 0.79 4.215 0.91 ;
        RECT 4.095 0.38 4.215 0.91 ;
        RECT 3.615 0.38 3.735 0.91 ;
        RECT 3.135 0.38 3.735 0.5 ;
        RECT 2.655 0.79 3.255 0.91 ;
        RECT 3.135 0.38 3.255 0.91 ;
        RECT 2.655 0.38 2.775 0.91 ;
        RECT 2.175 0.38 2.775 0.5 ;
        RECT 1.695 0.79 2.295 0.91 ;
        RECT 2.175 0.38 2.295 0.91 ;
        RECT 1.695 0.38 1.815 0.91 ;
        RECT 1.215 0.38 1.815 0.5 ;
        RECT 0.925 0.96 1.335 1.08 ;
        RECT 1.215 0.38 1.335 1.08 ;
        RECT 0.94 0.885 1.09 1.145 ;
        RECT 0.925 0.96 1.045 1.2 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.215 1.17 8.455 1.29 ;
        RECT 7.265 1.24 8.335 1.36 ;
        RECT 7.265 1.17 7.525 1.38 ;
        RECT 7.055 1.17 7.525 1.29 ;
    END
  END SN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7256 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.215 0.93 6.495 1.05 ;
        RECT 6.375 0.62 6.495 1.05 ;
        RECT 6.175 1.49 6.415 1.61 ;
        RECT 6.175 1.315 6.335 1.61 ;
        RECT 6.215 0.93 6.335 1.61 ;
        RECT 5.29 1.315 6.335 1.435 ;
        RECT 5.215 1.49 5.455 1.61 ;
        RECT 5.29 1.315 5.455 1.61 ;
        RECT 5.29 1.175 5.44 1.61 ;
        RECT 5.295 0.62 5.415 1.61 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.705 0.55 10.945 0.67 ;
        RECT 10.705 -0.18 10.825 0.67 ;
        RECT 8.415 0.45 8.655 0.57 ;
        RECT 8.535 -0.18 8.655 0.57 ;
        RECT 6.855 0.45 7.095 0.57 ;
        RECT 6.975 -0.18 7.095 0.57 ;
        RECT 5.775 0.45 6.015 0.57 ;
        RECT 5.895 -0.18 6.015 0.57 ;
        RECT 4.815 -0.18 4.935 0.67 ;
        RECT 3.855 -0.18 3.975 0.67 ;
        RECT 2.895 -0.18 3.015 0.67 ;
        RECT 1.935 -0.18 2.055 0.67 ;
        RECT 0.975 -0.18 1.095 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 10.925 1.795 11.045 2.79 ;
        RECT 9.295 2.23 9.535 2.79 ;
        RECT 8.515 2.23 8.635 2.79 ;
        RECT 7.675 2.23 7.795 2.79 ;
        RECT 6.655 1.98 6.895 2.1 ;
        RECT 6.655 1.98 6.775 2.79 ;
        RECT 5.695 1.97 5.935 2.09 ;
        RECT 5.695 1.97 5.815 2.79 ;
        RECT 4.735 1.97 4.975 2.09 ;
        RECT 4.735 1.97 4.855 2.79 ;
        RECT 3.775 1.97 4.015 2.09 ;
        RECT 3.775 1.97 3.895 2.79 ;
        RECT 2.815 1.97 3.055 2.09 ;
        RECT 2.815 1.97 2.935 2.79 ;
        RECT 1.855 1.97 2.095 2.09 ;
        RECT 1.855 1.97 1.975 2.79 ;
        RECT 0.955 2.07 1.075 2.79 ;
        RECT 0.135 1.55 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.465 1.915 11.345 1.915 11.345 0.91 10.31 0.91 10.31 0.81 10.045 0.81 10.045 0.48 9.925 0.48 9.925 0.36 10.165 0.36 10.165 0.69 10.43 0.69 10.43 0.79 11.245 0.79 11.245 0.62 11.365 0.62 11.365 0.74 11.465 0.74 ;
      POLYGON 11.205 1.675 10.645 1.675 10.645 2.155 10.045 2.155 10.045 2.11 7.71 2.11 7.71 1.86 6.385 1.86 6.385 1.85 0.555 1.85 0.555 1.5 0.685 1.5 0.685 0.98 0.275 0.98 0.275 0.62 0.395 0.62 0.395 0.86 0.805 0.86 0.805 1.73 6.505 1.73 6.505 1.74 7.83 1.74 7.83 1.99 10.045 1.99 10.045 1.63 9.545 1.63 9.545 1.17 9.665 1.17 9.665 1.51 10.165 1.51 10.165 2.035 10.525 2.035 10.525 1.15 10.145 1.15 10.145 1.03 10.645 1.03 10.645 1.555 11.085 1.555 11.085 1.335 11.205 1.335 ;
      POLYGON 10.405 1.915 10.285 1.915 10.285 1.39 9.905 1.39 9.905 1.05 8.095 1.05 8.095 1.12 7.855 1.12 7.855 0.93 9.705 0.93 9.705 0.62 9.825 0.62 9.825 0.93 10.025 0.93 10.025 1.27 10.405 1.27 ;
      RECT 8.815 1.75 9.925 1.87 ;
      POLYGON 9.215 1.43 8.695 1.43 8.695 1.62 8.155 1.62 8.155 1.87 8.035 1.87 8.035 1.62 6.815 1.62 6.815 1.29 6.455 1.29 6.455 1.17 6.815 1.17 6.815 0.93 7.615 0.93 7.615 0.62 7.735 0.62 7.735 1.05 6.935 1.05 6.935 1.5 8.035 1.5 8.035 1.48 8.155 1.48 8.155 1.5 8.575 1.5 8.575 1.31 9.215 1.31 ;
      POLYGON 4.495 1.61 4.255 1.61 4.255 1.49 4.335 1.49 4.335 1.15 3.495 1.15 3.495 1.49 3.535 1.49 3.535 1.61 3.295 1.61 3.295 1.49 3.375 1.49 3.375 1.15 2.655 1.15 2.655 1.03 3.375 1.03 3.375 0.62 3.495 0.62 3.495 1.03 4.335 1.03 4.335 0.62 4.455 0.62 4.455 1.49 4.495 1.49 ;
  END
END TLATSRX4

MACRO DFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX4 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.21 1.38 2.33 2.03 ;
        RECT 2.03 1.38 2.33 1.5 ;
        RECT 2.03 0.68 2.15 1.5 ;
        RECT 1.23 1.025 2.15 1.145 ;
        RECT 1.37 1.025 1.49 2.03 ;
        RECT 1.23 0.74 1.38 1.145 ;
        RECT 1.26 1.025 1.49 1.265 ;
        RECT 1.01 0.74 1.38 0.86 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.04 0.51 1.445 ;
        RECT 0.375 0.845 0.495 1.445 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.405 1.21 7.75 1.335 ;
        RECT 7.265 1.22 7.525 1.38 ;
    END
  END D
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.71 -0.18 7.83 0.83 ;
        RECT 5.71 0.49 5.95 0.61 ;
        RECT 5.83 -0.18 5.95 0.61 ;
        RECT 3.71 0.47 3.95 0.59 ;
        RECT 3.83 -0.18 3.95 0.59 ;
        RECT 2.51 0.47 2.75 0.59 ;
        RECT 2.51 -0.18 2.63 0.59 ;
        RECT 1.49 -0.18 1.73 0.32 ;
        RECT 0.53 -0.18 0.77 0.34 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.35 1.74 7.47 2.79 ;
        RECT 5.69 2.01 5.81 2.79 ;
        RECT 3.65 1.47 3.77 2.79 ;
        RECT 2.63 1.38 2.75 2.79 ;
        RECT 1.79 1.38 1.91 2.79 ;
        RECT 0.95 1.38 1.07 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.35 1.62 8.25 1.62 8.25 1.65 8.01 1.65 8.01 1.62 7.03 1.62 7.03 2.23 6.115 2.23 6.115 1.89 4.99 1.89 4.99 2.25 4.09 2.25 4.09 2.13 4.87 2.13 4.87 0.97 5.11 0.97 5.11 1.09 4.99 1.09 4.99 1.77 6.235 1.77 6.235 2.11 6.91 2.11 6.91 1.33 6.79 1.33 6.79 1.21 7.03 1.21 7.03 1.5 8.23 1.5 8.23 0.85 8.13 0.85 8.13 0.59 8.25 0.59 8.25 0.73 8.35 0.73 ;
      POLYGON 8.11 1.09 7.15 1.09 7.15 0.97 7.29 0.97 7.29 0.53 6.43 0.53 6.43 0.85 6.385 0.85 6.385 1.21 6.43 1.21 6.43 1.33 6.19 1.33 6.19 1.21 6.265 1.21 6.265 0.85 5.47 0.85 5.47 0.53 4.39 0.53 4.39 0.97 4.51 0.97 4.51 1.09 4.27 1.09 4.27 0.83 3.47 0.83 3.47 0.53 2.99 0.53 2.99 0.83 2.27 0.83 2.27 0.56 1.845 0.56 1.845 0.62 0.785 0.62 0.785 0.68 0.255 0.68 0.255 0.92 0.24 0.92 0.24 1.565 0.55 1.565 0.55 1.805 0.43 1.805 0.43 1.685 0.12 1.685 0.12 0.8 0.135 0.8 0.135 0.56 0.665 0.56 0.665 0.5 1.725 0.5 1.725 0.44 2.39 0.44 2.39 0.71 2.87 0.71 2.87 0.41 3.59 0.41 3.59 0.71 4.27 0.71 4.27 0.41 5.59 0.41 5.59 0.73 6.31 0.73 6.31 0.41 7.41 0.41 7.41 0.97 8.11 0.97 ;
      POLYGON 7.17 0.77 6.67 0.77 6.67 1.99 6.55 1.99 6.55 1.57 5.95 1.57 5.95 1.35 5.59 1.35 5.59 1.33 5.47 1.33 5.47 1.21 5.71 1.21 5.71 1.23 6.07 1.23 6.07 1.45 6.55 1.45 6.55 0.65 7.17 0.65 ;
      POLYGON 6.07 1.11 5.83 1.11 5.83 1.09 5.35 1.09 5.35 1.65 5.11 1.65 5.11 1.53 5.23 1.53 5.23 0.77 5.11 0.77 5.11 0.65 5.35 0.65 5.35 0.97 5.95 0.97 5.95 0.99 6.07 0.99 ;
      POLYGON 4.79 0.77 4.75 0.77 4.75 1.33 4.41 1.33 4.41 1.99 4.29 1.99 4.29 1.33 3.37 1.33 3.37 1.19 3.61 1.19 3.61 1.21 4.63 1.21 4.63 0.77 4.55 0.77 4.55 0.65 4.79 0.65 ;
      POLYGON 3.97 1.09 3.73 1.09 3.73 1.07 3.25 1.07 3.25 1.45 3.29 1.45 3.29 1.99 3.17 1.99 3.17 1.57 3.13 1.57 3.13 1.07 2.41 1.07 2.41 1.26 2.29 1.26 2.29 0.95 3.11 0.95 3.11 0.65 3.35 0.65 3.35 0.77 3.23 0.77 3.23 0.95 3.85 0.95 3.85 0.97 3.97 0.97 ;
  END
END DFFHQX4

MACRO AOI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X2 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 0.94 4.625 1.155 ;
        RECT 4.245 1.035 4.485 1.225 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.37 0.99 3.79 1.11 ;
        RECT 2.915 0.94 3.175 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.99 1.92 1.11 ;
        RECT 0.595 0.94 1.62 1.05 ;
        RECT 0.735 0.93 1.62 1.05 ;
        RECT 0.52 0.99 0.855 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.17 1.38 1.64 ;
        RECT 1.24 1.17 1.36 1.67 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.23 3.05 1.41 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6208 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 1.53 4.51 2.01 ;
        RECT 2.13 1.53 4.51 1.65 ;
        RECT 4.03 0.65 4.27 0.77 ;
        RECT 1.32 0.69 4.15 0.81 ;
        RECT 2.85 0.65 3.09 0.81 ;
        RECT 2.13 0.69 2.25 1.65 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.2 0.65 1.44 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 4.51 -0.18 4.63 0.64 ;
        RECT 3.55 0.45 3.79 0.57 ;
        RECT 3.55 -0.18 3.67 0.57 ;
        RECT 2.15 0.45 2.39 0.57 ;
        RECT 2.15 -0.18 2.27 0.57 ;
        RECT 0.62 -0.18 0.74 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 1.84 2.03 2.08 2.15 ;
        RECT 1.84 2.03 1.96 2.79 ;
        RECT 1 2.03 1.24 2.15 ;
        RECT 1 2.03 1.12 2.79 ;
        RECT 0.22 1.56 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.93 2.25 2.35 2.25 2.35 2.15 2.23 2.15 2.23 2.03 2.47 2.03 2.47 2.13 3.07 2.13 3.07 2.03 3.31 2.03 3.31 2.13 3.97 2.13 3.97 1.77 4.09 1.77 4.09 2.13 4.81 2.13 4.81 1.56 4.93 1.56 ;
      POLYGON 3.67 2.01 3.55 2.01 3.55 1.91 2.83 1.91 2.83 2.01 2.71 2.01 2.71 1.91 1.6 1.91 1.6 2.21 1.48 2.21 1.48 1.91 0.76 1.91 0.76 2.21 0.64 2.21 0.64 1.56 0.76 1.56 0.76 1.79 1.48 1.79 1.48 1.76 1.6 1.76 1.6 1.79 2.71 1.79 2.71 1.77 2.83 1.77 2.83 1.79 3.55 1.79 3.55 1.77 3.67 1.77 ;
  END
END AOI221X2

MACRO ADDFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX2 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4 0.83 6.515 0.95 ;
        RECT 3.125 0.76 4.12 0.88 ;
        RECT 3.205 0.65 3.465 0.88 ;
        RECT 3.125 0.71 3.245 0.95 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.975 1.07 7.235 1.38 ;
        RECT 2.875 1.07 7.235 1.19 ;
        RECT 3.815 1.07 4.055 1.2 ;
        RECT 1.865 1.02 2.995 1.14 ;
        RECT 1.745 1.08 1.985 1.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.64 1.31 6.855 1.43 ;
        RECT 2.635 1.32 4.88 1.44 ;
        RECT 3.55 1.32 3.7 1.725 ;
        RECT 3.275 1.31 3.555 1.44 ;
        RECT 2.165 1.26 2.755 1.38 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.68 0.765 2.21 ;
        RECT 0.36 1.175 0.765 1.295 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.695 0.885 8.05 1.145 ;
        RECT 7.635 1.62 7.875 2.15 ;
        RECT 7.695 0.64 7.815 2.15 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 8.115 -0.18 8.235 0.69 ;
        RECT 7.275 -0.18 7.395 0.69 ;
        RECT 5.065 0.35 5.305 0.47 ;
        RECT 5.065 -0.18 5.185 0.47 ;
        RECT 4.165 0.46 4.405 0.58 ;
        RECT 4.165 -0.18 4.285 0.58 ;
        RECT 1.965 -0.18 2.205 0.32 ;
        RECT 1.065 -0.18 1.185 0.73 ;
        RECT 0.225 -0.18 0.345 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 8.115 1.56 8.235 2.79 ;
        RECT 7.215 2.03 7.455 2.15 ;
        RECT 7.215 2.03 7.335 2.79 ;
        RECT 4.675 2.27 4.915 2.79 ;
        RECT 3.895 2.085 4.015 2.79 ;
        RECT 1.845 2 1.965 2.79 ;
        RECT 1.005 1.98 1.245 2.15 ;
        RECT 1.005 1.98 1.125 2.79 ;
        RECT 0.225 1.56 0.345 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.555 1.3 7.475 1.3 7.475 1.91 6.535 1.91 6.535 2.09 6.415 2.09 6.415 1.91 5.755 1.91 5.755 1.79 7.355 1.79 7.355 0.93 7.035 0.93 7.035 0.63 6.145 0.63 6.145 0.64 6.025 0.64 6.025 0.4 6.145 0.4 6.145 0.51 7.155 0.51 7.155 0.81 7.475 0.81 7.475 1.06 7.555 1.06 ;
      POLYGON 6.315 1.67 5.635 1.67 5.635 2.03 4.84 2.03 4.84 2.05 4.135 2.05 4.135 1.965 3.195 1.965 3.195 1.96 2.085 1.96 2.085 1.86 1.305 1.86 1.305 1.26 0.885 1.26 0.885 1.14 1.305 1.14 1.305 0.44 2.965 0.44 2.965 0.41 3.585 0.41 3.585 0.4 3.705 0.4 3.705 0.64 3.585 0.64 3.585 0.53 3.085 0.53 3.085 0.56 2.925 0.56 2.925 0.9 2.805 0.9 2.805 0.56 1.425 0.56 1.425 1.74 2.205 1.74 2.205 1.84 2.805 1.84 2.805 1.66 2.925 1.66 2.925 1.84 3.195 1.84 3.195 1.69 3.315 1.69 3.315 1.845 4.255 1.845 4.255 1.93 4.72 1.93 4.72 1.91 5.515 1.91 5.515 1.55 6.315 1.55 ;
      POLYGON 5.785 0.58 5.665 0.58 5.665 0.71 4.705 0.71 4.705 0.58 4.585 0.58 4.585 0.46 4.825 0.46 4.825 0.59 5.545 0.59 5.545 0.46 5.785 0.46 ;
      POLYGON 5.395 1.79 4.495 1.79 4.495 1.81 4.375 1.81 4.375 1.57 4.495 1.57 4.495 1.67 5.395 1.67 ;
      POLYGON 2.565 0.84 1.665 0.84 1.665 0.92 1.545 0.92 1.545 0.68 1.665 0.68 1.665 0.72 2.565 0.72 ;
      POLYGON 2.565 1.72 2.325 1.72 2.325 1.62 1.545 1.62 1.545 1.38 1.665 1.38 1.665 1.5 2.445 1.5 2.445 1.6 2.565 1.6 ;
  END
END ADDFX2

MACRO AOI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.68 0.82 1.04 ;
        RECT 0.65 0.5 0.8 0.855 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 0.5 1.38 0.96 ;
        RECT 1.21 0.47 1.33 0.96 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.57 0.8 1.69 1.235 ;
        RECT 1.52 0.885 1.67 1.3 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.785 0.51 1.24 ;
        RECT 0.36 0.76 0.48 1.24 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1932 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.48 1.515 1.72 ;
        RECT 1.215 1.48 1.515 1.6 ;
        RECT 1.215 1.08 1.335 1.6 ;
        RECT 0.97 1.08 1.335 1.2 ;
        RECT 0.94 0.885 1.09 1.145 ;
        RECT 0.97 0.4 1.09 1.2 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.71 -0.18 1.83 0.64 ;
        RECT 0.2 -0.18 0.32 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 0.555 1.6 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 1.84 1.755 1.84 1.755 1.96 0.975 1.96 0.975 1.48 0.315 1.48 0.315 1.66 0.075 1.66 0.075 1.54 0.195 1.54 0.195 1.36 1.095 1.36 1.095 1.84 1.635 1.84 1.635 1.72 1.815 1.72 1.815 1.6 1.935 1.6 ;
  END
END AOI22XL

MACRO TLATNTSCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX16 0 0 ;
  SIZE 14.21 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.845 0.565 1.1 ;
        RECT 0.265 0.98 0.505 1.21 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.76 1.09 1.205 ;
        RECT 0.925 0.76 1.045 1.23 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.76 1.385 1.25 ;
        RECT 1.23 0.76 1.385 1.22 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.535 1.345 13.655 2.205 ;
        RECT 8.48 1.225 13.555 1.345 ;
        RECT 13.435 0.655 13.555 1.465 ;
        RECT 12.655 0.775 13.555 0.895 ;
        RECT 12.695 1.225 12.815 2.205 ;
        RECT 12.535 0.725 12.775 0.845 ;
        RECT 11.855 1.225 11.975 2.205 ;
        RECT 11.755 0.655 11.875 1.345 ;
        RECT 10.975 0.775 11.875 0.895 ;
        RECT 11.015 1.225 11.135 2.21 ;
        RECT 10.855 0.725 11.095 0.845 ;
        RECT 10.175 1.225 10.295 2.21 ;
        RECT 10.075 0.655 10.195 1.345 ;
        RECT 9.295 0.775 10.195 0.895 ;
        RECT 9.335 1.225 9.455 2.21 ;
        RECT 9.175 0.725 9.415 0.845 ;
        RECT 8.48 1.175 8.63 1.435 ;
        RECT 8.495 0.785 8.615 2.21 ;
        RECT 8.395 0.665 8.515 0.905 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.21 0.18 ;
        RECT 13.855 -0.18 13.975 0.655 ;
        RECT 13.015 -0.18 13.135 0.655 ;
        RECT 12.175 -0.18 12.295 0.655 ;
        RECT 11.335 -0.18 11.455 0.655 ;
        RECT 10.495 -0.18 10.615 0.655 ;
        RECT 9.655 -0.18 9.775 0.655 ;
        RECT 8.815 -0.18 8.935 0.65 ;
        RECT 7.975 -0.18 8.095 0.65 ;
        RECT 6.455 0.47 6.695 0.59 ;
        RECT 6.455 -0.18 6.575 0.59 ;
        RECT 5.235 -0.18 5.355 0.76 ;
        RECT 4.155 -0.18 4.395 0.32 ;
        RECT 3.195 0.41 3.435 0.53 ;
        RECT 3.315 -0.18 3.435 0.53 ;
        RECT 1.005 -0.18 1.125 0.64 ;
        RECT 0.165 -0.18 0.285 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.21 2.79 ;
        RECT 13.955 1.465 14.075 2.79 ;
        RECT 13.115 1.465 13.235 2.79 ;
        RECT 12.275 1.465 12.395 2.79 ;
        RECT 11.435 1.465 11.555 2.79 ;
        RECT 10.595 1.465 10.715 2.79 ;
        RECT 9.755 1.465 9.875 2.79 ;
        RECT 8.915 1.465 9.035 2.79 ;
        RECT 8.075 1.72 8.195 2.79 ;
        RECT 7.235 1.72 7.355 2.79 ;
        RECT 6.395 1.72 6.515 2.79 ;
        RECT 5.555 1.72 5.675 2.79 ;
        RECT 4.715 1.69 4.835 2.79 ;
        RECT 3.815 2.23 3.935 2.79 ;
        RECT 2.765 1.98 3.005 2.1 ;
        RECT 2.765 1.98 2.885 2.79 ;
        RECT 0.885 1.61 1.005 2.79 ;
        RECT 0.765 1.61 1.005 1.73 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.275 1.24 8.135 1.24 8.135 1.6 7.775 1.6 7.775 2.21 7.655 2.21 7.655 1.6 6.935 1.6 6.935 2.21 6.815 2.21 6.815 1.6 6.095 1.6 6.095 2.21 5.975 2.21 5.975 1.6 5.255 1.6 5.255 2.21 5.135 2.21 5.135 1.48 8.015 1.48 8.015 1.12 7.375 1.12 7.375 0.84 7.235 0.84 7.235 0.83 5.935 0.83 5.935 0.78 5.815 0.78 5.815 0.66 6.055 0.66 6.055 0.71 7.235 0.71 7.235 0.6 7.355 0.6 7.355 0.72 7.495 0.72 7.495 1 8.275 1 ;
      POLYGON 7.895 1.36 4.595 1.36 4.595 1.81 4.415 1.81 4.415 2.21 4.295 2.21 4.295 1.69 4.475 1.69 4.475 1.31 3.155 1.31 3.155 1.37 3.035 1.37 3.035 1.13 3.155 1.13 3.155 1.19 4.635 1.19 4.635 0.68 4.875 0.68 4.875 0.8 4.755 0.8 4.755 1.24 7.895 1.24 ;
      POLYGON 7.255 1.12 5.575 1.12 5.575 1 4.995 1 4.995 0.56 4.515 0.56 4.515 0.64 4.035 0.64 4.035 0.76 3.915 0.76 3.915 1.01 2.915 1.01 2.915 1.49 3.485 1.49 3.485 1.75 3.605 1.75 3.605 1.87 3.365 1.87 3.365 1.61 2.795 1.61 2.795 1.26 2.715 1.26 2.715 0.89 3.795 0.89 3.795 0.64 3.915 0.64 3.915 0.52 4.395 0.52 4.395 0.44 5.115 0.44 5.115 0.88 5.695 0.88 5.695 1 7.255 1 ;
      POLYGON 4.355 1.55 4.175 1.55 4.175 2.11 3.125 2.11 3.125 1.86 2.645 1.86 2.645 1.92 2.305 1.92 2.305 2.04 2.185 2.04 2.185 1.92 2.105 1.92 2.105 0.74 2.235 0.74 2.235 0.62 2.355 0.62 2.355 0.86 2.225 0.86 2.225 1.8 2.525 1.8 2.525 1.74 3.245 1.74 3.245 1.99 4.055 1.99 4.055 1.43 4.355 1.43 ;
      POLYGON 3.795 0.48 3.675 0.48 3.675 0.77 2.955 0.77 2.955 0.5 2.595 0.5 2.595 1.1 2.465 1.1 2.465 1.62 2.345 1.62 2.345 0.98 2.475 0.98 2.475 0.5 1.625 0.5 1.625 1.61 1.365 1.61 1.365 1.49 1.505 1.49 1.505 0.64 1.425 0.64 1.425 0.38 2.035 0.38 2.035 0.36 2.275 0.36 2.275 0.38 3.075 0.38 3.075 0.65 3.555 0.65 3.555 0.36 3.795 0.36 ;
      POLYGON 1.935 1.94 1.885 1.94 1.885 2.06 1.765 2.06 1.765 1.94 1.125 1.94 1.125 1.49 0.305 1.49 0.305 1.67 0.185 1.67 0.185 1.37 0.685 1.37 0.685 0.725 0.585 0.725 0.585 0.4 0.705 0.4 0.705 0.605 0.805 0.605 0.805 1.37 1.245 1.37 1.245 1.82 1.815 1.82 1.815 0.62 1.935 0.62 ;
  END
END TLATNTSCAX16

MACRO NAND3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.765 0.99 2.885 1.42 ;
        RECT 2.68 1.025 2.83 1.44 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 2.025 0.99 2.22 1.23 ;
        RECT 0.805 0.99 2.22 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.23 1.435 1.5 ;
        RECT 1.125 1.23 1.435 1.48 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7616 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.56 2.405 2.21 ;
        RECT 0.305 1.62 2.405 1.74 ;
        RECT 1.445 1.62 1.565 2.21 ;
        RECT 0.305 0.51 1.525 0.63 ;
        RECT 0.605 1.56 0.725 2.21 ;
        RECT 0.305 1.56 0.725 1.74 ;
        RECT 0.305 1.52 0.565 1.74 ;
        RECT 0.305 0.51 0.425 1.74 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.445 0.46 2.685 0.58 ;
        RECT 2.445 -0.18 2.565 0.58 ;
        RECT 0.265 -0.18 0.505 0.39 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.705 1.56 2.825 2.79 ;
        RECT 1.865 1.86 1.985 2.79 ;
        RECT 1.025 1.86 1.145 2.79 ;
        RECT 0.185 1.86 0.305 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.305 1.8 3.185 1.8 3.185 1.68 3.005 1.68 3.005 0.87 2.56 0.87 2.56 1.17 2.44 1.17 2.44 0.87 0.665 0.87 0.665 1.17 0.545 1.17 0.545 0.75 2.985 0.75 2.985 0.59 3.105 0.59 3.105 0.71 3.125 0.71 3.125 1.56 3.305 1.56 ;
  END
END NAND3BX2

MACRO SDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRXL 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1.41 2.145 1.54 ;
        RECT 1.755 1.51 2.015 1.67 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.87 1.16 7.015 1.4 ;
        RECT 6.74 1.175 6.915 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.735 0.94 8.975 1.3 ;
        RECT 8.715 0.94 8.975 1.09 ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.155 0.94 9.555 1.17 ;
        RECT 9.155 0.94 9.275 1.35 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.675 0.96 10.135 1.15 ;
        RECT 9.875 0.935 10.135 1.15 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.405 1.32 1.525 1.91 ;
        RECT 1.365 0.68 1.485 0.96 ;
        RECT 1.23 1.175 1.445 1.435 ;
        RECT 1.325 0.84 1.445 1.44 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 9.015 -0.18 9.135 0.82 ;
        RECT 6.995 -0.18 7.115 0.84 ;
        RECT 4.945 -0.18 5.185 0.34 ;
        RECT 3.245 -0.18 3.485 0.34 ;
        RECT 1.785 -0.18 1.905 0.4 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 9.855 1.58 9.975 2.79 ;
        RECT 8.955 2.06 9.075 2.79 ;
        RECT 6.895 1.84 7.015 2.79 ;
        RECT 4.905 2.16 5.025 2.79 ;
        RECT 3.245 2.1 3.485 2.22 ;
        RECT 3.245 2.1 3.365 2.79 ;
        RECT 1.825 1.79 1.945 2.79 ;
        RECT 0.555 1.46 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.375 1.46 9.555 1.46 9.555 1.83 9.135 1.83 9.135 1.94 8.075 1.94 8.075 1.96 7.955 1.96 7.955 1.44 8.235 1.44 8.235 0.84 8.115 0.84 8.115 0.6 8.235 0.6 8.235 0.72 8.355 0.72 8.355 1.56 8.075 1.56 8.075 1.82 9.015 1.82 9.015 1.71 9.435 1.71 9.435 1.34 10.255 1.34 10.255 0.76 9.595 0.76 9.595 0.64 10.375 0.64 ;
      POLYGON 8.715 0.82 8.595 0.82 8.595 1.7 8.475 1.7 8.475 0.7 8.595 0.7 8.595 0.58 8.405 0.58 8.405 0.48 7.995 0.48 7.995 0.98 8.115 0.98 8.115 1.1 7.995 1.1 7.995 1.32 7.495 1.32 7.495 1.48 7.375 1.48 7.375 1.2 7.875 1.2 7.875 0.36 8.525 0.36 8.525 0.46 8.715 0.46 ;
      POLYGON 7.755 1.08 7.255 1.08 7.255 1.6 7.655 1.6 7.655 1.96 7.535 1.96 7.535 1.72 6.205 1.72 6.205 1.84 6.085 1.84 6.085 1.6 6.185 1.6 6.185 0.68 6.305 0.68 6.305 1.6 7.135 1.6 7.135 0.96 7.635 0.96 7.635 0.6 7.755 0.6 ;
      POLYGON 6.695 0.84 6.575 0.84 6.575 0.6 6.475 0.6 6.475 0.56 6.065 0.56 6.065 1.1 5.965 1.1 5.965 1.24 6.065 1.24 6.065 1.48 5.965 1.48 5.965 1.96 6.415 1.96 6.415 1.9 6.655 1.9 6.655 2.02 6.535 2.02 6.535 2.08 5.845 2.08 5.845 0.98 5.945 0.98 5.945 0.56 5.425 0.56 5.425 0.58 4.705 0.58 4.705 0.56 4.345 0.56 4.345 1.26 4.225 1.26 4.225 0.44 4.825 0.44 4.825 0.46 5.305 0.46 5.305 0.44 5.425 0.44 5.425 0.4 5.665 0.4 5.665 0.44 6.595 0.44 6.595 0.48 6.695 0.48 ;
      POLYGON 5.825 0.86 5.725 0.86 5.725 1.8 5.605 1.8 5.605 1.44 4.825 1.44 4.825 1.42 4.705 1.42 4.705 1.3 4.945 1.3 4.945 1.32 5.605 1.32 5.605 0.86 5.585 0.86 5.585 0.74 5.825 0.74 ;
      POLYGON 5.645 2.18 5.405 2.18 5.405 2.04 4.325 2.04 4.325 2.18 4.085 2.18 4.085 2.04 3.625 2.04 3.625 1.98 2.245 1.98 2.245 1.67 2.265 1.67 2.265 0.74 2.505 0.74 2.505 0.86 2.385 0.86 2.385 1.86 3.625 1.86 3.625 1.06 3.865 1.06 3.865 1.18 3.745 1.18 3.745 1.92 5.525 1.92 5.525 2.06 5.645 2.06 ;
      POLYGON 5.305 1.2 5.065 1.2 5.065 1.18 4.585 1.18 4.585 1.5 4.545 1.5 4.545 1.8 4.425 1.8 4.425 1.38 4.465 1.38 4.465 0.68 4.585 0.68 4.585 1.06 5.185 1.06 5.185 1.08 5.305 1.08 ;
      POLYGON 4.125 1.8 4.005 1.8 4.005 1.5 3.985 1.5 3.985 0.92 3.965 0.92 3.965 0.68 3.005 0.68 3.005 0.52 2.865 0.52 2.865 0.4 3.125 0.4 3.125 0.56 4.085 0.56 4.085 0.8 4.105 0.8 4.105 1.38 4.125 1.38 ;
      POLYGON 3.505 1.26 2.885 1.26 2.885 1.62 3.005 1.62 3.005 1.74 2.765 1.74 2.765 0.8 2.625 0.8 2.625 0.62 2.145 0.62 2.145 1.2 1.565 1.2 1.565 1.08 2.025 1.08 2.025 0.5 2.745 0.5 2.745 0.68 2.885 0.68 2.885 1.14 3.505 1.14 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END SDFFTRXL

MACRO OR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X2 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 0.51 1.455 ;
        RECT 0.375 1 0.495 1.485 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1.005 0.815 1.465 ;
        RECT 0.65 1 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.94 1.435 1.2 ;
        RECT 1.175 0.94 1.415 1.22 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.025 2.25 1.145 ;
        RECT 2.1 0.885 2.25 1.145 ;
        RECT 1.815 0.59 1.935 1.39 ;
        RECT 1.715 1.27 1.835 1.99 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 2.235 -0.18 2.355 0.64 ;
        RECT 1.335 0.46 1.575 0.58 ;
        RECT 1.335 -0.18 1.455 0.58 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 2.135 1.34 2.255 2.79 ;
        RECT 1.295 1.34 1.415 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.695 1.15 1.575 1.15 1.575 0.82 1.055 0.82 1.055 1.725 0.155 1.725 0.155 1.605 0.935 1.605 0.935 0.88 0.135 0.88 0.135 0.4 0.255 0.4 0.255 0.76 0.935 0.76 0.935 0.7 0.975 0.7 0.975 0.4 1.095 0.4 1.095 0.7 1.695 0.7 ;
  END
END OR3X2

MACRO CLKBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX2 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.225 1.275 1.38 ;
        RECT 1.155 1.13 1.275 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.225 0.675 2.12 ;
        RECT 0.555 0.605 0.675 0.845 ;
        RECT 0.515 0.725 0.635 1.345 ;
        RECT 0.36 0.885 0.635 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.77 ;
        RECT 0.135 -0.18 0.255 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.5 1.095 2.79 ;
        RECT 0.135 1.47 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.74 1.395 1.74 1.395 1.01 1.035 1.01 1.035 1.105 0.755 1.105 0.755 0.985 0.915 0.985 0.915 0.89 1.395 0.89 1.395 0.53 1.515 0.53 ;
  END
END CLKBUFX2

MACRO TLATX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX1 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.115 0.87 1.435 ;
        RECT 0.65 1.11 0.84 1.435 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1 3.41 1.47 ;
        RECT 3.26 1 3.38 1.5 ;
    END
  END G
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.94 0.59 4.06 2.21 ;
        RECT 3.84 0.885 4.06 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.17 0.68 5.29 2.12 ;
        RECT 4.945 0.94 5.29 1.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.75 -0.18 4.87 0.73 ;
        RECT 3.52 -0.18 3.64 0.64 ;
        RECT 2.23 -0.18 2.35 0.395 ;
        RECT 0.615 -0.18 0.735 0.395 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.75 1.47 4.87 2.79 ;
        RECT 3.52 1.62 3.64 2.79 ;
        RECT 1.93 2.215 2.17 2.79 ;
        RECT 0.59 1.795 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.05 1.33 4.45 1.33 4.45 2.12 4.33 2.12 4.33 0.68 4.45 0.68 4.45 1.21 5.05 1.21 ;
      POLYGON 3.72 1.22 3.6 1.22 3.6 0.88 2.83 0.88 2.83 1.515 2.65 1.515 2.65 1.855 2.41 1.855 2.41 1.735 2.53 1.735 2.53 1.515 1.93 1.515 1.93 1.395 2.71 1.395 2.71 0.675 2.83 0.675 2.83 0.76 3.72 0.76 ;
      POLYGON 3.22 0.64 3.1 0.64 3.1 0.555 2.59 0.555 2.59 0.635 1.94 0.635 1.94 0.615 1.43 0.615 1.43 1.475 1.21 1.475 1.21 1.595 1.11 1.595 1.11 2.075 1.52 2.075 1.52 1.975 3.04 1.975 3.04 1.68 3.16 1.68 3.16 2.095 1.64 2.095 1.64 2.195 0.99 2.195 0.99 1.675 0.41 1.675 0.41 1.335 0.53 1.335 0.53 1.555 0.99 1.555 0.99 1.355 1.31 1.355 1.31 0.495 1.71 0.495 1.71 0.395 1.95 0.395 1.95 0.495 2.06 0.495 2.06 0.515 2.47 0.515 2.47 0.435 3.1 0.435 3.1 0.4 3.22 0.4 ;
      POLYGON 2.49 1.275 1.67 1.275 1.67 1.835 1.35 1.835 1.35 1.955 1.23 1.955 1.23 1.715 1.55 1.715 1.55 0.735 1.79 0.735 1.79 0.855 1.67 0.855 1.67 1.155 2.49 1.155 ;
      POLYGON 1.19 1.235 1.07 1.235 1.07 0.99 0.29 0.99 0.29 1.915 0.17 1.915 0.17 0.915 0.135 0.915 0.135 0.675 0.255 0.675 0.255 0.795 0.29 0.795 0.29 0.87 1.19 0.87 ;
  END
END TLATX1

MACRO DFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX2 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1 0.405 1.24 ;
        RECT 0.07 1 0.405 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.12 1.755 1.355 ;
        RECT 1.175 1.12 1.435 1.38 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.515 0.64 5.635 1.18 ;
        RECT 5.455 1.06 5.575 2.21 ;
        RECT 5.29 1.175 5.575 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 5.995 -0.18 6.115 0.78 ;
        RECT 4.915 0.58 5.155 0.7 ;
        RECT 4.915 -0.18 5.035 0.7 ;
        RECT 3.015 0.58 3.255 0.7 ;
        RECT 3.015 -0.18 3.135 0.7 ;
        RECT 1.495 0.6 1.735 0.72 ;
        RECT 1.615 -0.18 1.735 0.72 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 5.875 1.56 5.995 2.79 ;
        RECT 5.035 1.56 5.155 2.79 ;
        RECT 3.215 2.23 3.455 2.79 ;
        RECT 1.415 1.76 1.535 2.79 ;
        RECT 0.145 1.46 0.265 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.535 1.44 6.475 1.44 6.475 2.08 6.355 2.08 6.355 1.44 5.755 1.44 5.755 1.2 5.875 1.2 5.875 1.32 6.415 1.32 6.415 0.64 6.535 0.64 ;
      POLYGON 6.235 1.2 6.115 1.2 6.115 1.02 5.755 1.02 5.755 0.52 5.395 0.52 5.395 0.94 4.895 0.94 4.895 1.42 4.615 1.42 4.615 1.81 4.455 1.81 4.455 2.21 4.335 2.21 4.335 1.69 4.495 1.69 4.495 1.3 4.775 1.3 4.775 0.94 4.66 0.94 4.66 0.8 4.275 0.8 4.275 0.68 4.78 0.68 4.78 0.82 5.275 0.82 5.275 0.4 5.875 0.4 5.875 0.9 6.235 0.9 ;
      POLYGON 4.655 1.18 3.975 1.18 3.975 1.61 3.855 1.61 3.855 1.06 3.875 1.06 3.875 0.5 3.495 0.5 3.495 0.94 2.855 0.94 2.855 1.59 2.735 1.59 2.735 0.56 2.015 0.56 2.015 0.96 2.035 0.96 2.035 1.4 1.915 1.4 1.915 1.08 1.895 1.08 1.895 0.96 1.255 0.96 1.255 0.56 0.685 0.56 0.685 1.58 0.565 1.58 0.565 0.44 1.155 0.44 1.155 0.36 1.395 0.36 1.395 0.48 1.375 0.48 1.375 0.84 1.895 0.84 1.895 0.44 2.855 0.44 2.855 0.82 3.375 0.82 3.375 0.38 3.995 0.38 3.995 1.06 4.655 1.06 ;
      POLYGON 4.375 1.57 4.215 1.57 4.215 2.11 2.905 2.11 2.905 2.25 2.255 2.25 2.255 1.64 1.055 1.64 1.055 2.09 0.935 2.09 0.935 0.8 0.895 0.8 0.895 0.68 1.135 0.68 1.135 0.8 1.055 0.8 1.055 1.52 2.255 1.52 2.255 1.35 2.375 1.35 2.375 2.13 2.785 2.13 2.785 1.99 4.095 1.99 4.095 1.45 4.255 1.45 4.255 1.33 4.375 1.33 ;
      POLYGON 3.935 1.87 3.615 1.87 3.615 1.19 3.015 1.19 3.015 1.07 3.615 1.07 3.615 0.74 3.635 0.74 3.635 0.62 3.755 0.62 3.755 0.86 3.735 0.86 3.735 1.75 3.935 1.75 ;
      POLYGON 3.495 1.83 2.615 1.83 2.615 2.01 2.495 2.01 2.495 0.8 2.135 0.8 2.135 0.68 2.615 0.68 2.615 1.71 3.375 1.71 3.375 1.35 3.495 1.35 ;
  END
END DFFHQX2

MACRO MXI4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4XL 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 0.48 2.455 1.08 ;
        RECT 2.315 0.96 2.435 1.47 ;
        RECT 0.68 0.48 2.455 0.6 ;
        RECT 1.835 0.4 2.075 0.6 ;
        RECT 0.68 1 0.84 1.24 ;
        RECT 0.68 0.48 0.8 1.24 ;
        RECT 0.65 0.595 0.8 0.855 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 1.26 3.275 1.46 ;
        RECT 2.915 1.155 3.175 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 1.51 4.535 1.65 ;
        RECT 4.075 1.5 4.335 1.67 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.655 1.44 4.915 1.67 ;
        RECT 4.695 1.26 4.815 1.67 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.955 1.55 6.235 1.7 ;
        RECT 5.815 1.5 6.075 1.685 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1752 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.9733 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.775 1.26 6.575 1.38 ;
        RECT 6.105 1.23 6.365 1.38 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.66 0.255 1.58 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.235 -0.18 6.355 0.38 ;
        RECT 4.555 -0.18 4.675 0.38 ;
        RECT 2.855 -0.18 2.975 0.86 ;
        RECT 1.31 -0.18 1.55 0.32 ;
        RECT 0.555 -0.18 0.795 0.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 6.135 1.96 6.255 2.79 ;
        RECT 4.685 2.03 4.805 2.79 ;
        RECT 4.565 2.03 4.805 2.15 ;
        RECT 2.895 2.14 3.015 2.79 ;
        RECT 1.255 1.91 1.375 2.79 ;
        RECT 1.135 1.91 1.375 2.03 ;
        RECT 0.555 2.04 0.795 2.16 ;
        RECT 0.555 2.04 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.825 0.9 6.815 0.9 6.815 1.62 6.675 1.62 6.675 2.08 6.555 2.08 6.555 1.5 6.695 1.5 6.695 0.78 6.705 0.78 6.705 0.62 5.995 0.62 5.995 0.54 5.415 0.54 5.415 1.67 5.295 1.67 5.295 0.62 4.31 0.62 4.31 0.56 3.635 0.56 3.635 1.54 3.395 1.54 3.395 1.42 3.515 1.42 3.515 0.44 3.935 0.44 3.935 0.36 4.175 0.36 4.175 0.44 4.43 0.44 4.43 0.5 5.295 0.5 5.295 0.42 5.615 0.42 5.615 0.4 5.855 0.4 5.855 0.42 6.115 0.42 6.115 0.5 6.825 0.5 ;
      POLYGON 5.655 1.96 5.575 1.96 5.575 2.08 5.455 2.08 5.455 1.96 4.925 1.96 4.925 1.91 4.25 1.91 4.25 2.25 3.335 2.25 3.335 2.13 3.135 2.13 3.135 2.02 2.675 2.02 2.675 2.25 2.555 2.25 2.555 1.9 3.255 1.9 3.255 2.01 3.455 2.01 3.455 2.13 4.13 2.13 4.13 1.79 5.045 1.79 5.045 1.84 5.535 1.84 5.535 0.66 5.655 0.66 ;
      POLYGON 5.175 1.16 4.935 1.16 4.935 1.14 4.115 1.14 4.115 1.38 3.995 1.38 3.995 1.02 5.175 1.02 ;
      POLYGON 4.035 0.8 3.875 0.8 3.875 1.89 3.715 1.89 3.715 2.01 3.595 2.01 3.595 1.89 3.375 1.89 3.375 1.78 2.435 1.78 2.435 2.11 1.735 2.11 1.735 2.25 1.495 2.25 1.495 2.13 1.615 2.13 1.615 1.99 2.315 1.99 2.315 1.66 3.495 1.66 3.495 1.77 3.755 1.77 3.755 0.68 4.035 0.68 ;
      POLYGON 2.215 0.84 2.195 0.84 2.195 1.75 2.175 1.75 2.175 1.87 2.055 1.87 2.055 1.76 0.38 1.76 0.38 1.02 0.5 1.02 0.5 1.64 2.055 1.64 2.055 1.63 2.075 1.63 2.075 0.84 1.975 0.84 1.975 0.72 2.215 0.72 ;
      POLYGON 1.955 1.47 1.225 1.47 1.225 1.52 0.985 1.52 0.985 1.4 1.04 1.4 1.04 0.84 0.92 0.84 0.92 0.72 1.16 0.72 1.16 1.35 1.835 1.35 1.835 1.23 1.955 1.23 ;
  END
END MXI4XL

MACRO AOI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X2 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.08 0.51 1.435 ;
        RECT 0.385 0.9 0.505 1.435 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.725 0.905 0.845 1.24 ;
        RECT 0.65 0.81 0.8 1.145 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.2 0.99 4.44 1.11 ;
        RECT 3.495 0.97 4.32 1.09 ;
        RECT 3.495 0.94 3.755 1.09 ;
        RECT 3.24 0.99 3.665 1.11 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.21 4.045 1.425 ;
        RECT 3.665 1.23 4.045 1.42 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.255 1.545 4.375 2.01 ;
        RECT 3 1.545 4.375 1.665 ;
        RECT 3.23 0.65 3.96 0.77 ;
        RECT 3.415 1.545 3.535 2.01 ;
        RECT 2.215 0.73 3.35 0.85 ;
        RECT 3 0.73 3.12 1.665 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 2.095 0.65 2.335 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.42 -0.18 4.54 0.64 ;
        RECT 2.87 0.46 3.11 0.58 ;
        RECT 2.87 -0.18 2.99 0.58 ;
        RECT 1.515 -0.18 1.635 0.64 ;
        RECT 0.555 -0.18 0.675 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 2.515 2.025 2.755 2.15 ;
        RECT 2.515 2.025 2.635 2.79 ;
        RECT 1.735 1.71 1.855 2.79 ;
        RECT 0.615 2.015 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.795 2.21 4.75 2.21 4.75 2.25 3.04 2.25 3.04 2.21 2.995 2.21 2.995 1.905 2.42 1.905 2.42 1.59 2.275 1.59 2.275 2.21 2.155 2.21 2.155 1.59 1.435 1.59 1.435 2.21 1.315 2.21 1.315 1.47 2.54 1.47 2.54 1.785 3.115 1.785 3.115 2.09 3.16 2.09 3.16 2.13 3.835 2.13 3.835 1.785 3.955 1.785 3.955 2.13 4.63 2.13 4.63 2.09 4.675 2.09 4.675 1.56 4.795 1.56 ;
      POLYGON 2.85 1.35 1.155 1.35 1.155 1.47 1.125 1.47 1.125 1.615 1.005 1.615 1.005 1.35 1.035 1.35 1.035 0.68 1.155 0.68 1.155 1.23 2.85 1.23 ;
      POLYGON 2.175 1.11 1.855 1.11 1.855 0.88 1.275 0.88 1.275 0.56 0.915 0.56 0.915 0.68 0.255 0.68 0.255 0.92 0.24 0.92 0.24 1.555 0.315 1.555 0.315 1.675 0.075 1.675 0.075 1.555 0.12 1.555 0.12 0.8 0.135 0.8 0.135 0.56 0.795 0.56 0.795 0.44 1.395 0.44 1.395 0.76 1.975 0.76 1.975 0.99 2.175 0.99 ;
  END
END AOI2BB2X2

MACRO NAND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X4 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.575 0.97 3.815 1.09 ;
        RECT 3.575 0.82 3.695 1.09 ;
        RECT 1.755 0.82 3.695 0.94 ;
        RECT 1.615 0.97 2.015 1.09 ;
        RECT 1.755 0.82 2.015 1.09 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.495 0.96 4.615 1.2 ;
        RECT 4.42 0.885 4.57 1.145 ;
        RECT 3.965 1.025 4.615 1.145 ;
        RECT 3.335 1.21 4.085 1.33 ;
        RECT 3.965 1.025 4.085 1.33 ;
        RECT 3.07 1.2 3.455 1.32 ;
        RECT 3.07 1.06 3.19 1.32 ;
        RECT 2.275 1.06 3.19 1.18 ;
        RECT 1.215 1.21 2.395 1.33 ;
        RECT 2.275 1.06 2.395 1.33 ;
        RECT 1.215 1.08 1.335 1.33 ;
        RECT 0.755 1.08 1.335 1.2 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.76 1.105 4.935 1.345 ;
        RECT 4.42 1.32 4.88 1.44 ;
        RECT 0.975 1.45 4.54 1.57 ;
        RECT 4.42 1.32 4.54 1.57 ;
        RECT 2.71 1.3 2.95 1.57 ;
        RECT 0.975 1.32 1.095 1.57 ;
        RECT 0.445 1.32 1.095 1.44 ;
        RECT 0.305 1.3 0.635 1.38 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.395 1.32 1.095 1.42 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.69 5.175 1.81 ;
        RECT 5.055 0.58 5.175 1.81 ;
        RECT 5 1.465 5.175 1.81 ;
        RECT 1.535 0.58 5.175 0.7 ;
        RECT 4.755 1.56 4.875 2.21 ;
        RECT 3.915 1.69 4.035 2.21 ;
        RECT 3.075 1.69 3.195 2.21 ;
        RECT 2.235 1.69 2.355 2.21 ;
        RECT 1.395 1.69 1.515 2.21 ;
        RECT 0.555 1.56 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.975 0.34 5.215 0.46 ;
        RECT 4.975 -0.18 5.095 0.46 ;
        RECT 2.555 0.34 2.795 0.46 ;
        RECT 2.555 -0.18 2.675 0.46 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 5.175 1.93 5.295 2.79 ;
        RECT 4.335 1.93 4.455 2.79 ;
        RECT 3.495 1.93 3.615 2.79 ;
        RECT 2.655 1.93 2.775 2.79 ;
        RECT 1.815 1.93 1.935 2.79 ;
        RECT 0.975 1.93 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND3X4

MACRO SDFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX2 0 0 ;
  SIZE 14.5 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.165 2.595 1.38 ;
        RECT 2.335 0.975 2.455 1.38 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.67 1.33 11.82 1.725 ;
        RECT 11.7 1.045 11.82 1.725 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.08 0.87 1.435 ;
        RECT 0.75 1.075 0.87 1.435 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.975 1.96 1.445 ;
        RECT 1.81 0.975 1.93 1.615 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7668 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.39 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.29 0.99 5.67 1.12 ;
        RECT 5.29 0.885 5.44 1.17 ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 0.755 1.21 0.995 ;
        RECT 0.94 0.595 1.09 0.955 ;
        RECT 0.37 0.835 1.21 0.955 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.4 0.68 12.52 2.205 ;
        RECT 12.25 1.465 12.52 1.725 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.24 1.545 13.48 1.665 ;
        RECT 13.3 0.68 13.42 1.085 ;
        RECT 13.24 0.965 13.36 1.665 ;
        RECT 13.065 1.23 13.36 1.38 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.5 0.18 ;
        RECT 13.72 -0.18 13.84 0.92 ;
        RECT 12.88 -0.18 13 0.73 ;
        RECT 11.86 -0.18 12.1 0.32 ;
        RECT 10.75 -0.18 10.87 0.78 ;
        RECT 6.03 -0.18 6.15 0.86 ;
        RECT 3.25 -0.18 3.49 0.74 ;
        RECT 2.05 0.495 2.29 0.615 ;
        RECT 2.17 -0.18 2.29 0.615 ;
        RECT 0.59 -0.18 0.71 0.675 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.5 2.79 ;
        RECT 13.72 2.025 13.96 2.145 ;
        RECT 13.72 2.025 13.84 2.79 ;
        RECT 12.76 2.025 13 2.145 ;
        RECT 12.76 2.025 12.88 2.79 ;
        RECT 11.98 1.845 12.1 2.79 ;
        RECT 10.81 2.2 10.93 2.79 ;
        RECT 9.29 1.94 9.41 2.79 ;
        RECT 6.89 1.98 7.13 2.13 ;
        RECT 6.89 1.98 7.01 2.79 ;
        RECT 5.57 1.8 5.69 2.79 ;
        RECT 3.3 1.72 3.54 1.84 ;
        RECT 3.3 1.72 3.42 2.79 ;
        RECT 1.87 1.735 1.99 2.79 ;
        RECT 0.53 2.23 0.65 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.32 2.085 14.2 2.085 14.2 1.325 13.5 1.325 13.5 1.205 14.14 1.205 14.14 0.68 14.26 0.68 14.26 1.205 14.32 1.205 ;
      POLYGON 14.08 1.905 12.825 1.905 12.825 1.455 12.64 1.455 12.64 0.56 12.28 0.56 12.28 1.26 12.16 1.26 12.16 0.56 11.29 0.56 11.29 0.68 11.31 0.68 11.31 1.52 11.29 1.52 11.29 1.84 11.17 1.84 11.17 1.4 11.19 1.4 11.19 1.02 10.21 1.02 10.21 1.1 10.09 1.1 10.09 0.86 10.21 0.86 10.21 0.9 11.17 0.9 11.17 0.44 12.76 0.44 12.76 1.215 12.945 1.215 12.945 1.785 13.96 1.785 13.96 1.505 14.08 1.505 ;
      POLYGON 11.68 0.925 11.55 0.925 11.55 1.845 11.68 1.845 11.68 2.085 11.56 2.085 11.56 2.08 10.79 2.08 10.79 1.82 10.115 1.82 10.115 2.01 9.77 2.01 9.77 1.89 9.995 1.89 9.995 1.7 10.91 1.7 10.91 1.96 11.43 1.96 11.43 0.805 11.56 0.805 11.56 0.68 11.68 0.68 ;
      POLYGON 11.07 1.26 10.95 1.26 10.95 1.34 8.45 1.34 8.45 1.72 8.33 1.72 8.33 0.68 8.57 0.68 8.57 0.8 8.45 0.8 8.45 1.22 10.83 1.22 10.83 1.14 11.07 1.14 ;
      POLYGON 10.67 2.06 10.55 2.06 10.55 2.25 9.53 2.25 9.53 1.82 9.17 1.82 9.17 1.9 8.905 1.9 8.905 1.96 8.45 1.96 8.45 2.14 7.25 2.14 7.25 1.86 6.77 1.86 6.77 2.25 5.89 2.25 5.89 2.13 6.65 2.13 6.65 1.74 7.37 1.74 7.37 2.02 8.33 2.02 8.33 1.84 8.785 1.84 8.785 1.78 9.05 1.78 9.05 1.7 9.65 1.7 9.65 2.13 10.43 2.13 10.43 1.94 10.67 1.94 ;
      POLYGON 10.51 1.58 8.93 1.58 8.93 1.66 8.69 1.66 8.69 1.54 8.81 1.54 8.81 1.46 10.51 1.46 ;
      POLYGON 10.45 0.78 10.33 0.78 10.33 0.54 10.21 0.54 10.21 0.48 9.73 0.48 9.73 0.54 9.61 0.54 9.61 0.78 9.49 0.78 9.49 0.42 9.61 0.42 9.61 0.36 10.33 0.36 10.33 0.42 10.45 0.42 ;
      POLYGON 10.09 0.72 9.97 0.72 9.97 1.02 8.81 1.02 8.81 0.62 8.93 0.62 8.93 0.9 9.85 0.9 9.85 0.6 10.09 0.6 ;
      POLYGON 8.71 0.48 8.21 0.48 8.21 1.9 7.49 1.9 7.49 1.62 6.53 1.62 6.53 2.01 5.81 2.01 5.81 1.68 5.24 1.68 5.24 2 5.09 2 5.09 2.2 4.85 2.2 4.85 2 3.78 2 3.78 1.64 3.87 1.64 3.87 0.86 3.85 0.86 3.85 0.74 4.09 0.74 4.09 0.86 3.99 0.86 3.99 1.76 3.9 1.76 3.9 1.88 4.47 1.88 4.47 1.4 4.49 1.4 4.49 0.98 4.61 0.98 4.61 1.52 4.59 1.52 4.59 1.88 5.12 1.88 5.12 1.56 5.93 1.56 5.93 1.89 6.41 1.89 6.41 1.5 7.61 1.5 7.61 1.78 8.09 1.78 8.09 0.36 8.71 0.36 ;
      POLYGON 7.97 1.66 7.73 1.66 7.73 1.54 7.85 1.54 7.85 1.38 6.17 1.38 6.17 1.65 6.29 1.65 6.29 1.77 6.05 1.77 6.05 1.44 5.21 1.44 5.21 1.32 6.05 1.32 6.05 1.26 6.87 1.26 6.87 0.62 6.99 0.62 6.99 1.26 7.85 1.26 7.85 0.62 7.97 0.62 ;
      POLYGON 7.41 0.86 7.29 0.86 7.29 0.5 6.75 0.5 6.75 0.62 6.57 0.62 6.57 0.86 6.45 0.86 6.45 0.5 6.63 0.5 6.63 0.38 7.41 0.38 ;
      POLYGON 6.69 1.14 5.79 1.14 5.79 0.765 4.95 0.765 4.95 1.76 4.71 1.76 4.71 1.64 4.83 1.64 4.83 0.8 4.71 0.8 4.71 0.68 4.83 0.68 4.83 0.645 5.91 0.645 5.91 1.02 6.69 1.02 ;
      POLYGON 4.45 0.86 4.35 0.86 4.35 1.76 4.11 1.76 4.11 1.64 4.23 1.64 4.23 0.74 4.33 0.74 4.33 0.62 3.73 0.62 3.73 0.98 3.01 0.98 3.01 0.495 2.53 0.495 2.53 0.855 1.81 0.855 1.81 0.635 1.45 0.635 1.45 1.915 1.17 1.915 1.17 1.795 1.33 1.795 1.33 0.435 1.45 0.435 1.45 0.515 1.93 0.515 1.93 0.735 2.41 0.735 2.41 0.375 3.13 0.375 3.13 0.86 3.61 0.86 3.61 0.5 4.45 0.5 ;
      POLYGON 3.75 1.22 2.89 1.22 2.89 1.795 2.23 1.795 2.23 1.675 2.77 1.675 2.77 0.735 2.65 0.735 2.65 0.615 2.89 0.615 2.89 1.1 3.75 1.1 ;
      POLYGON 1.69 2.155 0.93 2.155 0.93 1.675 0.255 1.675 0.255 1.83 0.135 1.83 0.135 1.71 0.13 1.71 0.13 0.595 0.17 0.595 0.17 0.435 0.29 0.435 0.29 0.715 0.25 0.715 0.25 1.555 1.09 1.555 1.09 1.295 1.21 1.295 1.21 1.675 1.05 1.675 1.05 2.035 1.57 2.035 1.57 0.755 1.69 0.755 ;
  END
END SDFFNSRX2

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 1.205 2.265 1.325 ;
        RECT 0.885 1.23 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.145 0.74 3.385 0.86 ;
        RECT 3.205 1.47 3.325 2.21 ;
        RECT 0.745 0.79 3.265 0.91 ;
        RECT 0.685 1.5 3.325 1.62 ;
        RECT 2.385 0.79 2.54 1.145 ;
        RECT 2.385 0.79 2.505 1.62 ;
        RECT 2.365 1.47 2.485 2.21 ;
        RECT 2.365 0.67 2.485 0.91 ;
        RECT 1.465 0.74 1.705 0.91 ;
        RECT 1.525 1.465 1.645 2.21 ;
        RECT 0.625 0.74 0.865 0.86 ;
        RECT 0.685 1.5 0.805 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.785 -0.18 2.905 0.67 ;
        RECT 1.945 -0.18 2.065 0.67 ;
        RECT 1.105 -0.18 1.225 0.67 ;
        RECT 0.265 -0.18 0.385 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.785 1.74 2.905 2.79 ;
        RECT 1.945 1.74 2.065 2.79 ;
        RECT 1.105 1.74 1.225 2.79 ;
        RECT 0.265 1.465 0.385 2.79 ;
    END
  END VDD
END INVX8

MACRO AOI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.57 1.03 1.69 1.455 ;
        RECT 1.52 1.03 1.69 1.435 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.885 1.09 1.185 ;
        RECT 0.85 0.88 0.97 1.17 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1 2.54 1.47 ;
        RECT 2.39 1 2.51 1.5 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.175 2.13 1.295 ;
        RECT 2.01 1.055 2.13 1.295 ;
        RECT 1.81 1.175 1.96 1.435 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1 1.38 1.455 ;
        RECT 1.23 1 1.35 1.485 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.76 0.51 1.235 ;
        RECT 0.36 0.76 0.51 1.215 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5276 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.465 2.83 1.725 ;
        RECT 2.69 1.465 2.81 2.21 ;
        RECT 2.68 0.76 2.8 1.74 ;
        RECT 1.85 1.62 2.81 1.74 ;
        RECT 1.43 0.76 2.8 0.88 ;
        RECT 1.85 1.56 1.97 2.01 ;
        RECT 1.43 0.59 1.55 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.49 -0.18 2.61 0.64 ;
        RECT 0.37 -0.18 0.49 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 1.01 1.845 1.13 2.79 ;
        RECT 0.17 1.56 0.29 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.39 2.25 1.43 2.25 1.43 1.725 0.71 1.725 0.71 2.21 0.59 2.21 0.59 1.56 0.71 1.56 0.71 1.605 1.55 1.605 1.55 2.13 2.27 2.13 2.27 1.86 2.39 1.86 ;
  END
END AOI33X1

MACRO OR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 1.025 1.96 1.145 ;
        RECT 1.81 0.885 1.96 1.145 ;
    END
  END A
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.03 0.51 1.485 ;
        RECT 0.36 1 0.48 1.485 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.05 0.82 1.485 ;
        RECT 0.7 1.025 0.82 1.485 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 1.105 1.155 1.46 ;
        RECT 0.94 1.135 1.09 1.485 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.075 0.59 3.195 0.83 ;
        RECT 2.055 1.505 3.175 1.625 ;
        RECT 3.075 0.59 3.175 1.625 ;
        RECT 2.895 1.505 3.12 1.725 ;
        RECT 2.97 1.465 3.175 1.625 ;
        RECT 3.055 0.71 3.12 1.725 ;
        RECT 2.235 0.76 3.175 0.88 ;
        RECT 2.895 1.505 3.015 2.21 ;
        RECT 2.235 0.59 2.355 0.88 ;
        RECT 2.055 1.505 2.175 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.495 -0.18 3.615 0.64 ;
        RECT 2.655 -0.18 2.775 0.64 ;
        RECT 1.815 -0.18 1.935 0.64 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.315 1.56 3.435 2.79 ;
        RECT 2.475 1.745 2.595 2.79 ;
        RECT 1.635 1.56 1.755 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.935 1.345 2.85 1.345 2.85 1.385 1.395 1.385 1.395 1.725 0.34 1.725 0.34 2.21 0.22 2.21 0.22 1.605 1.275 1.605 1.275 0.88 0.555 0.88 0.555 0.59 0.675 0.59 0.675 0.76 1.395 0.76 1.395 0.59 1.515 0.59 1.515 0.88 1.395 0.88 1.395 1.265 2.73 1.265 2.73 1.105 2.935 1.105 ;
  END
END OR4X4

MACRO DFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX1 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.905 1.21 2.145 1.44 ;
        RECT 1.755 1.23 2.015 1.485 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.795 2.13 7.675 2.25 ;
        RECT 6.795 1.78 6.915 2.25 ;
        RECT 5.595 1.78 6.915 1.9 ;
        RECT 5.115 1.84 5.715 1.96 ;
        RECT 5.115 1.7 5.235 1.96 ;
        RECT 4.005 1.7 5.235 1.82 ;
        RECT 3.255 1.77 4.125 1.89 ;
        RECT 3.255 1.52 3.465 1.89 ;
        RECT 3.255 1 3.375 1.89 ;
        RECT 3.205 1.52 3.465 1.67 ;
        RECT 3.135 1 3.375 1.12 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.435 0.835 9.79 1.21 ;
        RECT 9.435 0.835 9.555 1.22 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 0.865 10.66 1.32 ;
        RECT 10.52 0.865 10.64 1.34 ;
    END
  END CKN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 1.49 1.505 2.14 ;
        RECT 1.365 0.61 1.485 0.85 ;
        RECT 1.23 1.465 1.425 1.725 ;
        RECT 1.305 0.73 1.425 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.78 -0.18 10.9 0.745 ;
        RECT 9.43 -0.18 9.55 0.38 ;
        RECT 8.075 -0.18 8.315 0.36 ;
        RECT 3.075 -0.18 3.315 0.32 ;
        RECT 1.785 -0.18 1.905 0.85 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.78 1.46 10.9 2.79 ;
        RECT 9.355 1.9 9.475 2.79 ;
        RECT 7.815 2.13 7.935 2.79 ;
        RECT 6.075 2.26 6.315 2.79 ;
        RECT 4.485 2.18 4.725 2.3 ;
        RECT 4.485 2.18 4.605 2.79 ;
        RECT 3.165 2.25 3.405 2.79 ;
        RECT 1.805 1.605 1.925 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.48 0.745 10.39 0.745 10.39 1.46 10.48 1.46 10.48 1.7 10.36 1.7 10.36 1.58 10.27 1.58 10.27 0.6 9.79 0.6 9.79 0.62 9.14 0.62 9.14 0.6 7.635 0.6 7.635 0.48 7.515 0.48 7.515 0.36 7.755 0.36 7.755 0.48 8.615 0.48 8.615 0.38 8.855 0.38 8.855 0.48 9.26 0.48 9.26 0.5 9.67 0.5 9.67 0.38 9.99 0.38 9.99 0.48 10.48 0.48 ;
      POLYGON 10.15 0.84 10.03 0.84 10.03 1.46 9.915 1.46 9.915 2.02 9.795 2.02 9.795 1.46 9.135 1.46 9.135 2.2 8.415 2.2 8.415 2.01 7.035 2.01 7.035 1.66 6.715 1.66 6.715 1.44 6.305 1.44 6.305 1.32 6.835 1.32 6.835 1.54 7.155 1.54 7.155 1.89 8.535 1.89 8.535 2.08 9.015 2.08 9.015 1.46 8.675 1.46 8.675 1.53 8.555 1.53 8.555 1.29 8.675 1.29 8.675 1.34 9.015 1.34 9.015 1.28 9.275 1.28 9.275 1.34 9.91 1.34 9.91 0.72 10.15 0.72 ;
      POLYGON 9.015 0.84 8.895 0.84 8.895 1.17 8.435 1.17 8.435 1.65 8.775 1.65 8.775 1.84 8.895 1.84 8.895 1.96 8.655 1.96 8.655 1.77 8.315 1.77 8.315 1.17 7.195 1.17 7.195 1.05 8.775 1.05 8.775 0.72 9.015 0.72 ;
      POLYGON 8.195 1.56 7.955 1.56 7.955 1.42 7.395 1.42 7.395 1.65 7.515 1.65 7.515 1.77 7.275 1.77 7.275 1.42 6.955 1.42 6.955 1.14 6.185 1.14 6.185 1.66 5.845 1.66 5.845 1.54 6.065 1.54 6.065 0.86 5.945 0.86 5.945 0.62 6.065 0.62 6.065 0.74 6.185 0.74 6.185 1.02 6.955 1.02 6.955 0.78 7.035 0.78 7.035 0.66 7.155 0.66 7.155 0.9 7.075 0.9 7.075 1.3 8.075 1.3 8.075 1.44 8.195 1.44 ;
      POLYGON 7.635 0.84 7.395 0.84 7.395 0.72 7.275 0.72 7.275 0.54 6.865 0.54 6.865 0.66 6.735 0.66 6.735 0.9 6.615 0.9 6.615 0.54 6.745 0.54 6.745 0.42 7.395 0.42 7.395 0.6 7.515 0.6 7.515 0.72 7.635 0.72 ;
      POLYGON 6.675 2.23 6.435 2.23 6.435 2.14 5.955 2.14 5.955 2.2 4.875 2.2 4.875 2.06 4.365 2.06 4.365 2.13 4.345 2.13 4.345 2.25 4.225 2.25 4.225 2.13 2.655 2.13 2.655 2.085 2.225 2.085 2.225 1.725 2.265 1.725 2.265 0.61 2.385 0.61 2.385 1.845 2.345 1.845 2.345 1.965 2.775 1.965 2.775 2.01 4.245 2.01 4.245 1.94 4.995 1.94 4.995 2.08 5.835 2.08 5.835 2.02 6.555 2.02 6.555 2.11 6.675 2.11 ;
      POLYGON 5.945 1.34 5.705 1.34 5.705 0.48 5.265 0.48 5.265 0.36 5.825 0.36 5.825 1.22 5.945 1.22 ;
      POLYGON 5.585 0.86 5.475 0.86 5.475 1.72 5.355 1.72 5.355 1.34 3.495 1.34 3.495 0.88 3.015 0.88 3.015 1.24 3.035 1.24 3.035 1.36 2.795 1.36 2.795 1.24 2.895 1.24 2.895 0.76 3.615 0.76 3.615 1.22 5.355 1.22 5.355 0.74 5.465 0.74 5.465 0.62 5.585 0.62 ;
      POLYGON 5.165 1.1 4.235 1.1 4.235 0.62 4.355 0.62 4.355 0.98 5.045 0.98 5.045 0.62 5.165 0.62 ;
      POLYGON 5.115 1.58 3.885 1.58 3.885 1.65 3.645 1.65 3.645 1.53 3.765 1.53 3.765 1.46 5.115 1.46 ;
      POLYGON 4.775 0.86 4.655 0.86 4.655 0.5 4.115 0.5 4.115 0.72 3.975 0.72 3.975 0.8 3.735 0.8 3.735 0.68 3.855 0.68 3.855 0.6 3.995 0.6 3.995 0.38 4.775 0.38 ;
      POLYGON 3.875 0.48 3.735 0.48 3.735 0.56 2.775 0.56 2.775 0.86 2.675 0.86 2.675 1.52 2.865 1.52 2.865 1.76 2.745 1.76 2.745 1.64 2.555 1.64 2.555 0.74 2.655 0.74 2.655 0.56 2.555 0.56 2.555 0.49 2.145 0.49 2.145 1.09 1.785 1.09 1.785 1.11 1.545 1.11 1.545 0.97 2.025 0.97 2.025 0.37 2.675 0.37 2.675 0.44 3.615 0.44 3.615 0.36 3.875 0.36 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFNSRX1

MACRO NAND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.295 0.75 2.415 1.17 ;
        RECT 0.39 0.75 2.415 0.87 ;
        RECT 0.495 0.75 0.615 1.17 ;
        RECT 0.36 0.885 0.615 1.145 ;
        RECT 0.39 0.75 0.615 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.99 2.095 1.23 ;
        RECT 1.81 0.99 1.96 1.435 ;
        RECT 0.755 0.99 2.095 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.23 1.555 1.42 ;
        RECT 1.175 1.23 1.435 1.445 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7616 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.565 2.655 1.685 ;
        RECT 2.535 0.51 2.655 1.685 ;
        RECT 2.335 1.52 2.655 1.685 ;
        RECT 1.435 0.51 2.655 0.63 ;
        RECT 2.235 1.56 2.355 2.21 ;
        RECT 1.395 1.565 1.515 2.21 ;
        RECT 0.555 1.56 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.455 -0.18 2.695 0.39 ;
        RECT 0.275 0.46 0.515 0.58 ;
        RECT 0.275 -0.18 0.395 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.655 1.805 2.775 2.79 ;
        RECT 1.815 1.805 1.935 2.79 ;
        RECT 0.975 1.805 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND3X2

MACRO ADDFHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX4 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.035 0.82 7.495 0.94 ;
        RECT 5.175 0.82 5.415 1.09 ;
        RECT 4.055 0.78 5.155 0.9 ;
        RECT 4.075 0.65 4.335 0.9 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 0.94 8.395 1.25 ;
        RECT 8.135 0.94 8.395 1.16 ;
        RECT 7.655 1.04 8.395 1.16 ;
        RECT 5.535 1.06 7.775 1.18 ;
        RECT 4.795 1.21 5.655 1.33 ;
        RECT 5.535 1.06 5.655 1.33 ;
        RECT 4.795 1.02 4.915 1.33 ;
        RECT 3.735 1.02 4.915 1.14 ;
        RECT 2.675 0.98 3.855 1.1 ;
        RECT 2.675 0.98 2.795 1.24 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.895 1.28 8.135 1.4 ;
        RECT 5.775 1.3 8.015 1.42 ;
        RECT 4.42 1.45 5.895 1.57 ;
        RECT 5.775 1.3 5.895 1.57 ;
        RECT 4.42 1.28 4.675 1.57 ;
        RECT 4.42 1.28 4.57 1.725 ;
        RECT 4.05 1.28 4.675 1.4 ;
        RECT 3.135 1.26 4.17 1.34 ;
        RECT 3.255 1.28 4.675 1.38 ;
        RECT 3.135 1.22 3.375 1.34 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.32 1.555 2.21 ;
        RECT 1.435 0.67 1.555 0.96 ;
        RECT 0.555 1.32 1.555 1.44 ;
        RECT 0.555 0.84 1.555 0.96 ;
        RECT 0.595 1.32 0.715 2.21 ;
        RECT 0.595 0.67 0.715 0.96 ;
        RECT 0.555 0.79 0.675 1.44 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.735 0.885 10.08 1.145 ;
        RECT 8.855 1.32 9.855 1.44 ;
        RECT 9.735 0.76 9.855 1.44 ;
        RECT 9.695 1.32 9.815 2.21 ;
        RECT 8.855 0.76 9.855 0.88 ;
        RECT 9.695 0.59 9.815 0.88 ;
        RECT 8.855 1.32 8.975 2.21 ;
        RECT 8.855 0.59 8.975 0.88 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 10.115 -0.18 10.235 0.64 ;
        RECT 9.275 -0.18 9.395 0.64 ;
        RECT 8.375 0.46 8.615 0.58 ;
        RECT 8.375 -0.18 8.495 0.58 ;
        RECT 5.935 0.34 6.175 0.46 ;
        RECT 5.935 -0.18 6.055 0.46 ;
        RECT 5.095 -0.18 5.215 0.64 ;
        RECT 2.815 -0.18 3.055 0.38 ;
        RECT 1.855 -0.18 1.975 0.72 ;
        RECT 1.015 -0.18 1.135 0.72 ;
        RECT 0.175 -0.18 0.295 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 10.115 1.56 10.235 2.79 ;
        RECT 9.275 1.56 9.395 2.79 ;
        RECT 8.375 2.02 8.615 2.15 ;
        RECT 8.375 2.02 8.495 2.79 ;
        RECT 5.935 2.17 6.175 2.79 ;
        RECT 4.975 2.17 5.215 2.79 ;
        RECT 2.875 2.1 2.995 2.79 ;
        RECT 1.795 2.03 2.035 2.15 ;
        RECT 1.795 2.03 1.915 2.79 ;
        RECT 1.015 1.56 1.135 2.79 ;
        RECT 0.175 1.56 0.295 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.615 1.12 8.635 1.12 8.635 1.9 7.655 1.9 7.655 2.15 7.415 2.15 7.415 1.9 7.255 1.9 7.255 2.15 7.015 2.15 7.015 1.88 7.135 1.88 7.135 1.78 8.515 1.78 8.515 0.82 8.135 0.82 8.135 0.7 6.835 0.7 6.835 0.58 7.515 0.58 7.515 0.5 7.755 0.5 7.755 0.58 8.255 0.58 8.255 0.7 8.635 0.7 8.635 1 9.615 1 ;
      POLYGON 7.335 1.66 6.895 1.66 6.895 2.05 4.455 2.05 4.455 2.21 4.335 2.21 4.335 2.05 3.895 2.05 3.895 2.15 3.775 2.15 3.775 2.05 3.685 2.05 3.685 1.98 2.36 1.98 2.36 1.91 2.095 1.91 2.095 1.2 0.795 1.2 0.795 1.08 2.095 1.08 2.095 0.5 3.775 0.5 3.775 0.41 4.575 0.41 4.575 0.65 4.455 0.65 4.455 0.53 3.895 0.53 3.895 0.74 3.775 0.74 3.775 0.62 2.215 0.62 2.215 1.79 2.48 1.79 2.48 1.86 3.775 1.86 3.775 1.5 3.895 1.5 3.895 1.93 4.335 1.93 4.335 1.845 4.455 1.845 4.455 1.93 6.775 1.93 6.775 1.54 7.335 1.54 ;
      RECT 5.455 0.58 6.655 0.7 ;
      POLYGON 6.655 1.81 5.455 1.81 5.455 1.69 6.415 1.69 6.415 1.62 6.655 1.62 ;
      RECT 2.335 0.74 3.535 0.86 ;
      POLYGON 3.475 1.74 3.355 1.74 3.355 1.62 2.515 1.62 2.515 1.67 2.395 1.67 2.395 1.34 2.515 1.34 2.515 1.5 3.475 1.5 ;
  END
END ADDFHX4

MACRO SEDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX2 0 0 ;
  SIZE 14.79 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.39 1.98 1.41 ;
        RECT 0.9 0.39 1.98 0.51 ;
        RECT 0.3 0.97 1.22 1.09 ;
        RECT 0.9 0.39 1.02 1.09 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.23 0.88 1.47 ;
        RECT 0.595 1.21 0.855 1.47 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.32 1.175 7.47 1.585 ;
        RECT 7.35 1.1 7.47 1.585 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.23 10.735 1.48 ;
        RECT 10.455 1.23 10.715 1.5 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.745 1.18 13.865 1.42 ;
        RECT 12.75 1.26 13.865 1.38 ;
        RECT 13.355 1.23 13.615 1.38 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.225 1.15 14.485 1.42 ;
        RECT 14.225 1.02 14.465 1.42 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.09 1.175 8.34 1.435 ;
        RECT 8.07 0.74 8.31 0.86 ;
        RECT 8.09 0.74 8.21 1.48 ;
        RECT 8.04 1.36 8.16 1.68 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9 0.74 9.27 0.86 ;
        RECT 9 0.74 9.12 1.68 ;
        RECT 8.77 1.175 9.12 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.79 0.18 ;
        RECT 14.115 -0.18 14.235 0.82 ;
        RECT 12.43 0.51 12.67 0.63 ;
        RECT 12.43 -0.18 12.55 0.63 ;
        RECT 12.1 -0.18 12.22 0.63 ;
        RECT 10.86 -0.18 11.1 0.32 ;
        RECT 9.51 -0.18 9.75 0.38 ;
        RECT 8.55 -0.18 8.79 0.38 ;
        RECT 7.59 -0.18 7.83 0.34 ;
        RECT 6.24 0.53 6.48 0.65 ;
        RECT 6.24 -0.18 6.36 0.65 ;
        RECT 4.24 0.55 4.48 0.67 ;
        RECT 4.36 -0.18 4.48 0.67 ;
        RECT 2.14 -0.18 2.26 0.81 ;
        RECT 0.56 -0.18 0.68 0.81 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.79 2.79 ;
        RECT 14.055 2.16 14.175 2.79 ;
        RECT 10.875 2.01 10.995 2.79 ;
        RECT 10.755 2.01 10.995 2.13 ;
        RECT 9.48 2.08 9.6 2.79 ;
        RECT 8.46 2.04 8.7 2.16 ;
        RECT 8.46 2.04 8.58 2.79 ;
        RECT 7.56 2.21 7.68 2.79 ;
        RECT 6.17 2.29 6.41 2.79 ;
        RECT 4.01 2.23 4.13 2.79 ;
        RECT 2.34 2.29 2.58 2.79 ;
        RECT 0.62 1.83 0.86 1.95 ;
        RECT 0.62 1.83 0.74 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.725 1.66 14.655 1.66 14.655 1.9 14.14 1.9 14.14 2.04 13.61 2.04 13.61 2.18 13.105 2.18 13.105 2.06 13.49 2.06 13.49 1.92 14.02 1.92 14.02 1.78 14.535 1.78 14.535 1.54 14.605 1.54 14.605 0.9 14.535 0.9 14.535 0.58 14.655 0.58 14.655 0.78 14.725 0.78 ;
      POLYGON 14.105 1.66 13.815 1.66 13.815 1.78 13.695 1.78 13.695 1.54 13.985 1.54 13.985 1.06 13.695 1.06 13.695 0.48 12.91 0.48 12.91 0.87 12.035 0.87 12.035 1.26 11.915 1.26 11.915 0.75 12.79 0.75 12.79 0.36 13.815 0.36 13.815 0.94 14.105 0.94 ;
      POLYGON 13.425 1.8 13.305 1.8 13.305 1.62 12.63 1.62 12.63 1.68 12.585 1.68 12.585 1.8 12.465 1.8 12.465 1.5 10.975 1.5 10.975 1.89 10.635 1.89 10.635 2.25 9.72 2.25 9.72 1.92 7.455 1.92 7.455 2.09 6.05 2.09 6.05 2.25 4.25 2.25 4.25 2.11 3.89 2.11 3.89 2.17 2.14 2.17 2.14 2.15 2.02 2.15 2.02 2.03 2.26 2.03 2.26 2.05 3.77 2.05 3.77 1.99 4.37 1.99 4.37 2.13 5.93 2.13 5.93 1.97 7.335 1.97 7.335 1.8 9.84 1.8 9.84 2.13 10.515 2.13 10.515 1.77 10.855 1.77 10.855 1.38 11.46 1.38 11.46 0.86 11.34 0.86 11.34 0.74 11.58 0.74 11.58 1.38 12.51 1.38 12.51 0.99 13.13 0.99 13.13 0.6 13.37 0.6 13.37 0.72 13.25 0.72 13.25 1.11 12.63 1.11 12.63 1.5 13.425 1.5 ;
      POLYGON 13.065 1.86 12.945 1.86 12.945 2.04 12.57 2.04 12.57 2.25 11.655 2.25 11.655 1.95 11.775 1.95 11.775 2.13 12.45 2.13 12.45 1.92 12.825 1.92 12.825 1.74 13.065 1.74 ;
      POLYGON 12.255 2.01 12.015 2.01 12.015 1.83 11.535 1.83 11.535 2.01 11.175 2.01 11.175 1.89 11.415 1.89 11.415 1.71 12.135 1.71 12.135 1.89 12.255 1.89 ;
      POLYGON 11.74 0.52 11.395 0.52 11.395 0.56 10.07 0.56 10.07 0.62 7.95 0.62 7.95 0.98 7.97 0.98 7.97 1.24 7.85 1.24 7.85 1.1 7.83 1.1 7.83 0.62 6.9 0.62 6.9 0.86 6.79 0.86 6.79 1.49 6.87 1.49 6.87 1.61 6.63 1.61 6.63 1.45 5.93 1.45 5.93 1.33 6.67 1.33 6.67 0.74 6.78 0.74 6.78 0.5 9.87 0.5 9.87 0.4 10.11 0.4 10.11 0.44 11.275 0.44 11.275 0.4 11.74 0.4 ;
      POLYGON 11.135 1.18 10.855 1.18 10.855 1.11 10.335 1.11 10.335 1.89 10.395 1.89 10.395 2.01 10.155 2.01 10.155 1.89 10.215 1.89 10.215 0.98 10.44 0.98 10.44 0.68 10.56 0.68 10.56 0.99 10.975 0.99 10.975 1.06 11.135 1.06 ;
      POLYGON 10.23 0.86 10.095 0.86 10.095 1.3 10.025 1.3 10.025 1.68 9.905 1.68 9.905 1.3 9.24 1.3 9.24 1.18 9.975 1.18 9.975 0.74 10.23 0.74 ;
      POLYGON 7.35 0.86 7.2 0.86 7.2 1.85 5.81 1.85 5.81 2.01 4.49 2.01 4.49 1.69 3.81 1.69 3.81 1.27 3.93 1.27 3.93 1.57 4.61 1.57 4.61 1.89 5.09 1.89 5.09 1.45 5.07 1.45 5.07 1.33 5.31 1.33 5.31 1.45 5.21 1.45 5.21 1.89 5.69 1.89 5.69 1.13 5.68 1.13 5.68 1.01 5.92 1.01 5.92 1.13 5.81 1.13 5.81 1.73 7.08 1.73 7.08 0.74 7.35 0.74 ;
      POLYGON 6.55 1.2 6.43 1.2 6.43 0.89 5.56 0.89 5.56 1.65 5.57 1.65 5.57 1.77 5.33 1.77 5.33 1.65 5.44 1.65 5.44 0.74 5.48 0.74 5.48 0.62 5.6 0.62 5.6 0.74 5.755 0.74 5.755 0.77 6.55 0.77 ;
      POLYGON 5.32 1.18 5.2 1.18 5.2 0.56 4.72 0.56 4.72 0.91 4 0.91 4 0.5 3.42 0.5 3.42 1.51 3.3 1.51 3.3 0.5 2.89 0.5 2.89 0.57 2.68 0.57 2.68 0.69 2.74 0.69 2.74 1.57 2.94 1.57 2.94 1.69 2.62 1.69 2.62 0.81 2.56 0.81 2.56 0.45 2.77 0.45 2.77 0.38 3.68 0.38 3.68 0.36 3.92 0.36 3.92 0.38 4.12 0.38 4.12 0.79 4.6 0.79 4.6 0.44 5.32 0.44 ;
      POLYGON 5.08 1.15 4.95 1.15 4.95 1.65 4.97 1.65 4.97 1.77 4.73 1.77 4.73 1.65 4.83 1.65 4.83 1.45 4.11 1.45 4.11 1.33 4.83 1.33 4.83 1.03 4.84 1.03 4.84 0.68 5.08 0.68 ;
      POLYGON 4.71 1.15 3.69 1.15 3.69 1.83 3.57 1.83 3.57 0.8 3.54 0.8 3.54 0.68 3.78 0.68 3.78 0.8 3.69 0.8 3.69 1.03 4.71 1.03 ;
      POLYGON 3.27 1.93 2.38 1.93 2.38 1.91 1.6 1.91 1.6 1.55 1.62 1.55 1.62 0.75 1.14 0.75 1.14 0.63 1.74 0.63 1.74 1.67 1.72 1.67 1.72 1.79 2.5 1.79 2.5 1.81 3.06 1.81 3.06 0.62 3.18 0.62 3.18 1.63 3.27 1.63 ;
      POLYGON 1.5 1.43 1.48 1.43 1.48 1.71 0.32 1.71 0.32 1.83 0.2 1.83 0.2 1.71 0.06 1.71 0.06 0.69 0.14 0.69 0.14 0.57 0.26 0.57 0.26 0.81 0.18 0.81 0.18 1.59 1.36 1.59 1.36 1.31 1.38 1.31 1.38 1.19 1.5 1.19 ;
  END
END SEDFFTRX2

MACRO NOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X8 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.855 1.05 5.095 1.17 ;
        RECT 0.68 0.965 4.975 1.085 ;
        RECT 3.495 0.965 3.735 1.17 ;
        RECT 1.995 0.965 2.235 1.17 ;
        RECT 0.65 1.055 0.8 1.435 ;
        RECT 0.435 1.055 0.8 1.175 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.375 1.19 5.835 1.31 ;
        RECT 1.315 1.29 5.495 1.41 ;
        RECT 5.235 1.23 5.835 1.31 ;
        RECT 3.995 1.21 4.235 1.41 ;
        RECT 2.735 1.205 2.975 1.41 ;
        RECT 1.195 1.205 1.435 1.325 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.53 6.075 1.65 ;
        RECT 5.955 0.71 6.075 1.65 ;
        RECT 5.815 1.47 6.02 1.725 ;
        RECT 5.87 1.465 6.075 1.65 ;
        RECT 0.495 0.71 6.075 0.83 ;
        RECT 5.815 1.47 5.935 2.21 ;
        RECT 4.335 1.53 4.455 2.21 ;
        RECT 2.535 1.53 2.655 2.21 ;
        RECT 1.175 1.53 1.295 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.955 0.46 6.195 0.58 ;
        RECT 5.955 -0.18 6.075 0.58 ;
        RECT 5.115 0.46 5.355 0.58 ;
        RECT 5.115 -0.18 5.235 0.58 ;
        RECT 4.275 0.46 4.515 0.58 ;
        RECT 4.275 -0.18 4.395 0.58 ;
        RECT 3.435 0.46 3.675 0.58 ;
        RECT 3.435 -0.18 3.555 0.58 ;
        RECT 2.595 0.46 2.835 0.58 ;
        RECT 2.595 -0.18 2.715 0.58 ;
        RECT 1.755 0.46 1.995 0.58 ;
        RECT 1.755 -0.18 1.875 0.58 ;
        RECT 0.915 0.46 1.155 0.58 ;
        RECT 0.915 -0.18 1.035 0.58 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.175 1.77 5.295 2.79 ;
        RECT 3.295 1.77 3.415 2.79 ;
        RECT 1.895 1.77 2.015 2.79 ;
        RECT 0.335 1.465 0.455 2.79 ;
    END
  END VDD
END NOR2X8

MACRO AOI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32XL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.775 0.51 1.235 ;
        RECT 0.38 0.775 0.5 1.265 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.175 0.995 2.295 1.435 ;
        RECT 2.1 0.775 2.25 1.195 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 0.725 1.16 1.055 ;
        RECT 0.94 0.595 1.09 0.93 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.655 0.615 1.775 1.055 ;
        RECT 1.52 0.775 1.67 1.195 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.735 0.82 1.105 ;
        RECT 0.65 0.49 0.8 0.855 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2388 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.315 2.055 1.675 ;
        RECT 1.23 1.315 2.055 1.435 ;
        RECT 1.32 0.415 1.44 0.655 ;
        RECT 1.23 1.175 1.4 1.435 ;
        RECT 1.28 0.535 1.4 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 2.155 -0.18 2.275 0.655 ;
        RECT 0.22 -0.18 0.34 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.095 2.075 1.215 2.79 ;
        RECT 0.135 2.075 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.475 1.795 2.295 1.795 2.295 1.915 1.515 1.915 1.515 1.675 0.555 1.675 0.555 1.555 1.635 1.555 1.635 1.795 2.175 1.795 2.175 1.675 2.355 1.675 2.355 1.555 2.475 1.555 ;
  END
END AOI32XL

MACRO OAI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X4 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.055 1.06 7.175 1.18 ;
        RECT 4.13 1.06 4.28 1.435 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.535 0.99 3.695 1.11 ;
        RECT 2.915 0.94 3.175 1.11 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.675 1.3 6.195 1.42 ;
        RECT 4.655 1.52 4.915 1.67 ;
        RECT 4.675 1.3 4.915 1.67 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 1.26 3.035 1.38 ;
        RECT 2.625 1.23 2.885 1.38 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.855 0.65 7.095 0.77 ;
        RECT 4.335 0.76 6.975 0.88 ;
        RECT 6.015 0.65 6.255 0.88 ;
        RECT 5.875 1.56 5.995 2.21 ;
        RECT 1.735 1.79 5.995 1.91 ;
        RECT 5.175 0.65 5.415 0.88 ;
        RECT 4.595 1.79 4.715 2.21 ;
        RECT 4.335 0.65 4.575 0.88 ;
        RECT 3.815 0.82 4.455 0.94 ;
        RECT 3.785 1.79 4.045 1.96 ;
        RECT 3.815 0.82 3.935 1.96 ;
        RECT 3.115 1.56 3.235 2.21 ;
        RECT 1.735 1.56 1.855 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 3.435 0.34 3.675 0.46 ;
        RECT 3.435 -0.18 3.555 0.46 ;
        RECT 2.475 0.34 2.715 0.46 ;
        RECT 2.475 -0.18 2.595 0.46 ;
        RECT 1.515 0.34 1.755 0.46 ;
        RECT 1.515 -0.18 1.635 0.46 ;
        RECT 0.555 0.34 0.795 0.46 ;
        RECT 0.555 -0.18 0.675 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.515 1.56 6.635 2.79 ;
        RECT 5.175 2.03 5.415 2.15 ;
        RECT 5.175 2.03 5.295 2.79 ;
        RECT 3.795 2.08 4.035 2.2 ;
        RECT 3.795 2.08 3.915 2.79 ;
        RECT 2.315 2.03 2.555 2.15 ;
        RECT 2.315 2.03 2.435 2.79 ;
        RECT 1.095 1.56 1.215 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.455 0.65 7.335 0.65 7.335 0.53 6.615 0.53 6.615 0.64 6.495 0.64 6.495 0.53 5.775 0.53 5.775 0.64 5.655 0.64 5.655 0.53 4.935 0.53 4.935 0.64 4.815 0.64 4.815 0.53 4.095 0.53 4.095 0.7 0.075 0.7 0.075 0.58 3.975 0.58 3.975 0.41 4.815 0.41 4.815 0.4 4.935 0.4 4.935 0.41 5.655 0.41 5.655 0.4 5.775 0.4 5.775 0.41 6.495 0.41 6.495 0.4 6.615 0.4 6.615 0.41 7.455 0.41 ;
  END
END OAI22X4

MACRO NOR4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBXL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.12 0.565 1.38 ;
        RECT 0.305 1.04 0.545 1.38 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.23 2.885 1.445 ;
        RECT 2.505 1.325 2.745 1.515 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.615 1.265 1.735 1.55 ;
        RECT 1.52 1.43 1.67 1.725 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.995 1.24 1.115 1.665 ;
        RECT 0.94 1.315 1.09 1.725 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2544 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.075 1.175 2.25 1.435 ;
        RECT 2.095 0.4 2.215 0.64 ;
        RECT 1.075 1.845 2.195 1.965 ;
        RECT 2.075 0.52 2.195 1.965 ;
        RECT 1.255 0.76 2.195 0.88 ;
        RECT 1.255 0.4 1.375 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.515 -0.18 2.635 0.64 ;
        RECT 1.675 -0.18 1.795 0.64 ;
        RECT 0.775 -0.18 0.895 0.53 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.315 1.84 2.435 2.79 ;
        RECT 0.135 1.5 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.125 1.9 2.675 1.9 2.675 1.78 3.005 1.78 3.005 0.98 2.315 0.98 2.315 0.86 3.005 0.86 3.005 0.64 2.935 0.64 2.935 0.4 3.055 0.4 3.055 0.52 3.125 0.52 ;
      POLYGON 1.955 1.12 0.805 1.12 0.805 1.62 0.675 1.62 0.675 1.74 0.555 1.74 0.555 1.5 0.685 1.5 0.685 0.92 0.525 0.92 0.525 0.68 0.645 0.68 0.645 0.8 0.805 0.8 0.805 1 1.955 1 ;
  END
END NOR4BBXL

MACRO SDFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX4 0 0 ;
  SIZE 14.5 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.445 1.515 2.095 ;
        RECT 1.395 0.63 1.515 0.97 ;
        RECT 1.375 0.85 1.495 1.565 ;
        RECT 0.555 0.97 1.495 1.09 ;
        RECT 0.555 0.94 0.855 1.09 ;
        RECT 0.555 0.63 0.675 2.095 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.005 3.12 1.455 ;
        RECT 2.97 0.98 3.09 1.455 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.43 1.265 11.55 1.515 ;
        RECT 11.035 1.265 11.55 1.385 ;
        RECT 11.035 1.23 11.295 1.385 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.67 1.28 12.015 1.485 ;
        RECT 11.67 1.09 11.82 1.485 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.315 1.235 13.615 1.465 ;
        RECT 13.355 1.21 13.615 1.465 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.985 0.97 14.105 1.22 ;
        RECT 12.735 0.97 14.105 1.09 ;
        RECT 13.645 0.94 13.905 1.09 ;
        RECT 12.735 0.97 12.975 1.1 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 2.13 8.555 2.25 ;
        RECT 7.675 2.01 8.435 2.13 ;
        RECT 7.675 1.7 7.795 2.13 ;
        RECT 7.075 1.7 7.795 1.82 ;
        RECT 5.755 2.13 7.195 2.25 ;
        RECT 7.075 1.7 7.195 2.25 ;
        RECT 5.755 1.52 5.875 2.25 ;
        RECT 5.235 1.52 5.875 1.64 ;
        RECT 5.235 1.52 5.495 1.67 ;
        RECT 5.055 1.47 5.355 1.59 ;
    END
  END SN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.5 0.18 ;
        RECT 14.245 -0.18 14.365 0.88 ;
        RECT 13.235 0.46 13.475 0.58 ;
        RECT 13.235 -0.18 13.355 0.58 ;
        RECT 11.815 -0.18 12.055 0.34 ;
        RECT 11.185 -0.18 11.425 0.38 ;
        RECT 9.135 0.46 9.375 0.58 ;
        RECT 9.135 -0.18 9.255 0.58 ;
        RECT 5.205 -0.18 5.325 0.46 ;
        RECT 2.595 0.5 2.835 0.62 ;
        RECT 2.715 -0.18 2.835 0.62 ;
        RECT 1.815 -0.18 1.935 0.68 ;
        RECT 0.975 -0.18 1.095 0.68 ;
        RECT 0.135 -0.18 0.255 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.5 2.79 ;
        RECT 14.245 1.46 14.365 2.79 ;
        RECT 13.515 1.825 13.635 2.79 ;
        RECT 12.235 1.76 12.355 2.79 ;
        RECT 10.975 1.94 11.095 2.79 ;
        RECT 8.675 2.01 8.915 2.13 ;
        RECT 8.675 2.01 8.795 2.79 ;
        RECT 7.315 1.94 7.555 2.06 ;
        RECT 7.315 1.94 7.435 2.79 ;
        RECT 4.855 2.29 5.095 2.79 ;
        RECT 3.595 2.175 3.715 2.79 ;
        RECT 2.715 2.175 2.835 2.79 ;
        RECT 1.815 1.575 1.935 2.79 ;
        RECT 0.975 1.445 1.095 2.79 ;
        RECT 0.135 1.445 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.005 0.82 13.355 0.82 13.355 0.85 12.615 0.85 12.615 1.22 13.135 1.22 13.135 1.585 13.765 1.585 13.765 1.495 14.005 1.495 14.005 1.615 13.885 1.615 13.885 1.705 13.015 1.705 13.015 1.34 12.495 1.34 12.495 1.1 12.375 1.1 12.375 0.98 12.495 0.98 12.495 0.73 13.235 0.73 13.235 0.7 14.005 0.7 ;
      POLYGON 12.995 2.21 12.875 2.21 12.875 1.945 12.775 1.945 12.775 1.58 12.135 1.58 12.135 0.61 11.725 0.61 11.725 0.62 10.945 0.62 10.945 0.48 10.375 0.48 10.375 0.72 10.195 0.72 10.195 1.8 10.175 1.8 10.175 2.01 10.055 2.01 10.055 1.68 10.075 1.68 10.075 0.36 11.065 0.36 11.065 0.5 11.605 0.5 11.605 0.49 12.755 0.49 12.755 0.61 12.255 0.61 12.255 1.46 12.895 1.46 12.895 1.825 12.995 1.825 ;
      POLYGON 11.995 1.94 11.49 1.94 11.49 1.82 10.65 1.82 10.65 2.25 9.395 2.25 9.395 1.89 7.915 1.89 7.915 1.58 6.955 1.58 6.955 2.01 6.235 2.01 6.235 1.29 6.275 1.29 6.275 0.91 6.355 0.91 6.355 0.55 5.875 0.55 5.875 1.11 5.635 1.11 5.635 0.99 5.755 0.99 5.755 0.43 6.475 0.43 6.475 1.03 6.395 1.03 6.395 1.41 6.355 1.41 6.355 1.89 6.835 1.89 6.835 1.46 8.035 1.46 8.035 1.77 9.395 1.77 9.395 1.42 9.675 1.42 9.675 1.54 9.515 1.54 9.515 2.13 10.53 2.13 10.53 1.7 10.795 1.7 10.795 1.1 10.775 1.1 10.775 0.86 11.43 0.86 11.43 0.74 11.695 0.74 11.695 0.86 11.55 0.86 11.55 0.98 10.915 0.98 10.915 1.7 11.61 1.7 11.61 1.82 11.995 1.82 ;
      POLYGON 10.825 0.72 10.615 0.72 10.615 1.46 10.675 1.46 10.675 1.58 10.435 1.58 10.435 1.46 10.495 1.46 10.495 1.32 10.315 1.32 10.315 1.08 10.495 1.08 10.495 0.6 10.825 0.6 ;
      POLYGON 9.955 0.74 9.935 0.74 9.935 1.78 9.755 1.78 9.755 2.01 9.635 2.01 9.635 1.66 9.815 1.66 9.815 0.74 9.69 0.74 9.69 0.82 8.875 0.82 8.875 1 8.635 1 8.635 0.88 8.755 0.88 8.755 0.7 9.57 0.7 9.57 0.62 9.835 0.62 9.835 0.5 9.955 0.5 ;
      POLYGON 9.695 1.24 8.395 1.24 8.395 1.1 6.835 1.1 6.835 0.98 8.515 0.98 8.515 1.12 9.455 1.12 9.455 1.1 9.695 1.1 ;
      POLYGON 9.275 1.54 8.415 1.54 8.415 1.65 8.155 1.65 8.155 1.34 6.715 1.34 6.715 1.77 6.475 1.77 6.475 1.53 6.595 1.53 6.595 0.6 6.715 0.6 6.715 0.74 7.955 0.74 7.955 0.6 8.195 0.6 8.195 0.72 8.075 0.72 8.075 0.86 6.715 0.86 6.715 1.22 8.275 1.22 8.275 1.42 9.275 1.42 ;
      POLYGON 8.555 0.68 8.435 0.68 8.435 0.48 7.835 0.48 7.835 0.62 7.535 0.62 7.535 0.5 7.715 0.5 7.715 0.36 8.555 0.36 ;
      POLYGON 6.235 0.79 6.115 0.79 6.115 1.99 5.995 1.99 5.995 1.35 4.815 1.35 4.815 1.57 4.315 1.57 4.315 2.01 3.695 2.01 3.695 2.055 2.515 2.055 2.515 1.255 2.635 1.255 2.635 1.935 3.575 1.935 3.575 1.89 4.195 1.89 4.195 1.45 4.695 1.45 4.695 1.23 5.995 1.23 5.995 0.67 6.235 0.67 ;
      POLYGON 5.635 0.79 5.395 0.79 5.395 0.7 4.965 0.7 4.965 0.48 4.485 0.48 4.485 0.5 4.425 0.5 4.425 0.62 4.185 0.62 4.185 0.5 4.305 0.5 4.305 0.38 4.365 0.38 4.365 0.36 5.085 0.36 5.085 0.58 5.515 0.58 5.515 0.67 5.635 0.67 ;
      POLYGON 5.635 1.93 4.435 1.93 4.435 1.69 4.555 1.69 4.555 1.81 5.395 1.81 5.395 1.79 5.635 1.79 ;
      POLYGON 5.635 2.25 5.215 2.25 5.215 2.17 4.645 2.17 4.645 2.25 3.875 2.25 3.875 2.13 4.525 2.13 4.525 2.05 5.335 2.05 5.335 2.13 5.635 2.13 ;
      POLYGON 4.845 0.86 4.575 0.86 4.575 1.28 3.705 1.28 3.705 0.72 3.585 0.72 3.585 0.6 3.825 0.6 3.825 1.16 4.455 1.16 4.455 0.74 4.605 0.74 4.605 0.6 4.845 0.6 ;
      POLYGON 4.335 1.04 4.095 1.04 4.095 0.86 3.945 0.86 3.945 0.48 3.075 0.48 3.075 0.86 2.355 0.86 2.355 2.095 2.235 2.095 2.235 1.21 1.615 1.21 1.615 1.09 2.235 1.09 2.235 0.54 2.355 0.54 2.355 0.74 2.955 0.74 2.955 0.36 4.065 0.36 4.065 0.74 4.215 0.74 4.215 0.92 4.335 0.92 ;
      POLYGON 3.585 1.33 3.36 1.33 3.36 1.695 3.315 1.695 3.315 1.815 3.195 1.815 3.195 1.575 3.24 1.575 3.24 0.72 3.195 0.72 3.195 0.6 3.435 0.6 3.435 0.72 3.36 0.72 3.36 1.21 3.585 1.21 ;
  END
END SDFFSRHQX4

MACRO TBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX20 0 0 ;
  SIZE 19.72 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.08 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.085 0.94 10.865 1.06 ;
        RECT 6.085 0.76 6.205 1.06 ;
        RECT 5.665 0.76 6.205 0.88 ;
        RECT 5.665 0.41 5.785 0.88 ;
        RECT 5.065 0.41 5.785 0.53 ;
        RECT 4.585 0.785 5.185 0.905 ;
        RECT 5.065 0.41 5.185 0.905 ;
        RECT 4.865 0.785 4.985 1.15 ;
        RECT 4.585 0.36 4.705 0.905 ;
        RECT 3.885 0.36 4.705 0.48 ;
        RECT 2.945 0.78 4.005 0.9 ;
        RECT 3.885 0.36 4.005 0.9 ;
        RECT 3.385 0.78 3.505 1.1 ;
        RECT 2.945 0.36 3.065 0.9 ;
        RECT 2.085 0.36 3.065 0.48 ;
        RECT 1.605 0.78 2.205 0.9 ;
        RECT 2.085 0.36 2.205 0.9 ;
        RECT 2.025 0.78 2.145 1.12 ;
        RECT 1.625 0.78 1.745 1.12 ;
        RECT 1.605 0.36 1.725 0.9 ;
        RECT 0.605 0.36 1.725 0.48 ;
        RECT 0.305 0.94 0.725 1.06 ;
        RECT 0.605 0.36 0.725 1.06 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3926 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.756 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.5193 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.845 1.22 4.225 1.34 ;
        RECT 4.105 1.07 4.225 1.34 ;
        RECT 2.915 1.22 3.175 1.38 ;
        RECT 2.845 1.07 2.965 1.34 ;
    END
  END OE
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 19.045 1.4 19.165 2.17 ;
        RECT 17.245 0.76 19.045 0.88 ;
        RECT 18.925 0.59 19.045 0.88 ;
        RECT 18.865 1.4 19.165 1.52 ;
        RECT 11.665 1.28 18.985 1.4 ;
        RECT 18.865 0.76 18.985 1.52 ;
        RECT 18.205 1.28 18.325 2.17 ;
        RECT 18.085 0.59 18.205 0.88 ;
        RECT 17.365 1.28 17.485 2.17 ;
        RECT 17.245 0.59 17.365 0.88 ;
        RECT 16.525 1.28 16.645 2.17 ;
        RECT 16.405 0.59 16.525 1.4 ;
        RECT 15.565 0.76 16.525 0.88 ;
        RECT 15.685 1.28 15.805 2.17 ;
        RECT 15.565 0.59 15.685 0.88 ;
        RECT 14.845 1.28 14.965 2.17 ;
        RECT 14.725 0.59 14.845 0.83 ;
        RECT 14.545 0.71 14.845 0.83 ;
        RECT 14.545 0.71 14.665 1.4 ;
        RECT 13.885 0.76 14.665 0.88 ;
        RECT 14.005 1.28 14.125 2.17 ;
        RECT 13.885 0.59 14.005 0.88 ;
        RECT 13.165 1.28 13.285 2.17 ;
        RECT 13.045 0.59 13.165 0.83 ;
        RECT 12.865 0.71 13.165 0.83 ;
        RECT 12.865 0.71 12.985 1.4 ;
        RECT 12.205 0.76 12.985 0.88 ;
        RECT 12.325 1.28 12.445 2.17 ;
        RECT 12.205 0.59 12.325 0.88 ;
        RECT 11.67 0.885 11.82 1.145 ;
        RECT 11.665 0.92 11.79 1.4 ;
        RECT 11.485 1.52 11.785 1.64 ;
        RECT 11.665 0.92 11.785 1.64 ;
        RECT 11.365 0.92 11.82 1.04 ;
        RECT 11.485 1.52 11.605 2.17 ;
        RECT 11.365 0.59 11.485 1.04 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 19.72 0.18 ;
        RECT 19.345 -0.18 19.465 0.64 ;
        RECT 18.505 -0.18 18.625 0.64 ;
        RECT 17.665 -0.18 17.785 0.64 ;
        RECT 16.825 -0.18 16.945 0.64 ;
        RECT 15.985 -0.18 16.105 0.64 ;
        RECT 15.145 -0.18 15.265 0.64 ;
        RECT 14.305 -0.18 14.425 0.64 ;
        RECT 13.465 -0.18 13.585 0.64 ;
        RECT 12.625 -0.18 12.745 0.64 ;
        RECT 11.785 -0.18 11.905 0.64 ;
        RECT 10.885 0.46 11.125 0.58 ;
        RECT 10.885 -0.18 11.005 0.58 ;
        RECT 10.045 0.46 10.285 0.58 ;
        RECT 10.045 -0.18 10.165 0.58 ;
        RECT 9.205 0.46 9.445 0.58 ;
        RECT 9.205 -0.18 9.325 0.58 ;
        RECT 8.365 0.46 8.605 0.58 ;
        RECT 8.365 -0.18 8.485 0.58 ;
        RECT 7.525 0.46 7.765 0.58 ;
        RECT 7.525 -0.18 7.645 0.58 ;
        RECT 6.685 0.46 6.925 0.58 ;
        RECT 6.685 -0.18 6.805 0.58 ;
        RECT 5.905 -0.18 6.025 0.64 ;
        RECT 4.825 -0.18 4.945 0.665 ;
        RECT 3.325 -0.18 3.445 0.66 ;
        RECT 1.845 -0.18 1.965 0.66 ;
        RECT 0.365 -0.18 0.485 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 19.72 2.79 ;
        RECT 19.465 1.52 19.585 2.79 ;
        RECT 18.625 1.52 18.745 2.79 ;
        RECT 17.785 1.52 17.905 2.79 ;
        RECT 16.945 1.52 17.065 2.79 ;
        RECT 16.105 1.52 16.225 2.79 ;
        RECT 15.265 1.52 15.385 2.79 ;
        RECT 14.425 1.52 14.545 2.79 ;
        RECT 13.585 1.52 13.705 2.79 ;
        RECT 12.745 1.52 12.865 2.79 ;
        RECT 11.905 1.52 12.025 2.79 ;
        RECT 11.005 1.9 11.245 2.11 ;
        RECT 11.005 1.9 11.125 2.79 ;
        RECT 9.165 1.9 9.405 2.02 ;
        RECT 9.165 1.9 9.285 2.79 ;
        RECT 7.505 2.055 7.745 2.175 ;
        RECT 7.505 2.055 7.625 2.79 ;
        RECT 6.105 2.01 6.345 2.13 ;
        RECT 6.105 2.01 6.225 2.79 ;
        RECT 5.205 1.51 5.325 2.79 ;
        RECT 4.305 2.23 4.425 2.79 ;
        RECT 3.585 2.23 3.705 2.79 ;
        RECT 2.745 2.23 2.865 2.79 ;
        RECT 1.905 2.23 2.025 2.79 ;
        RECT 1.065 2.23 1.185 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.445 1.4 11.365 1.4 11.365 1.78 10.57 1.78 10.57 2.25 9.525 2.25 9.525 1.78 9.045 1.78 9.045 2.25 7.865 2.25 7.865 1.935 6.54 1.935 6.54 1.89 5.445 1.89 5.445 1.39 4.905 1.39 4.905 1.95 4.785 1.95 4.785 1.62 4.065 1.62 4.065 1.95 3.945 1.95 3.945 1.62 3.225 1.62 3.225 1.95 3.105 1.95 3.105 1.62 2.385 1.62 2.385 1.95 2.265 1.95 2.265 1.62 1.545 1.62 1.545 1.95 1.425 1.95 1.425 1.62 0.705 1.62 0.705 1.95 0.585 1.95 0.585 1.405 0.705 1.405 0.705 1.5 0.945 1.5 0.945 0.6 1.185 0.6 1.185 0.72 1.065 0.72 1.065 1.5 1.425 1.5 1.425 1.48 1.545 1.48 1.545 1.5 2.265 1.5 2.265 1.48 2.385 1.48 2.385 1.5 2.605 1.5 2.605 0.72 2.585 0.72 2.585 0.6 2.825 0.6 2.825 0.72 2.725 0.72 2.725 1.5 3.945 1.5 3.945 1.46 4.065 1.46 4.065 1.5 4.345 1.5 4.345 0.72 4.125 0.72 4.125 0.6 4.465 0.6 4.465 1.5 4.785 1.5 4.785 1.27 5.565 1.27 5.565 1.77 6.66 1.77 6.66 1.815 7.985 1.815 7.985 2.13 8.925 2.13 8.925 1.66 9.645 1.66 9.645 2.13 10.45 2.13 10.45 1.66 11.245 1.66 11.245 1.28 11.325 1.28 11.325 1.16 11.445 1.16 ;
      POLYGON 11.125 1.17 11.105 1.17 11.105 1.54 10.225 1.54 10.225 2.01 10.105 2.01 10.105 1.54 8.545 1.54 8.545 2.01 8.425 2.01 8.425 1.54 7.045 1.54 7.045 1.695 6.805 1.695 6.805 1.575 6.925 1.575 6.925 1.42 10.985 1.42 10.985 0.82 6.325 0.82 6.325 0.52 6.445 0.52 6.445 0.7 7.165 0.7 7.165 0.52 7.285 0.52 7.285 0.7 8.005 0.7 8.005 0.52 8.125 0.52 8.125 0.7 8.845 0.7 8.845 0.52 8.965 0.52 8.965 0.7 9.685 0.7 9.685 0.515 9.805 0.515 9.805 0.7 10.525 0.7 10.525 0.515 10.645 0.515 10.645 0.7 11.105 0.7 11.105 0.93 11.125 0.93 ;
      POLYGON 10.005 1.3 5.805 1.3 5.805 1.65 5.685 1.65 5.685 1.12 5.305 1.12 5.305 0.65 5.545 0.65 5.545 1 5.805 1 5.805 1.18 10.005 1.18 ;
      POLYGON 2.485 1.36 1.285 1.36 1.285 1.085 1.405 1.085 1.405 1.24 2.365 1.24 2.365 1.09 2.485 1.09 ;
  END
END TBUFX20

MACRO INVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX16 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.728 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.205 5.495 1.325 ;
        RECT 0.885 1.205 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.5 5.735 1.62 ;
        RECT 5.615 0.79 5.735 1.62 ;
        RECT 5.58 1.465 5.73 1.725 ;
        RECT 5.595 1.465 5.715 2.21 ;
        RECT 0.615 0.79 5.735 0.91 ;
        RECT 5.595 0.67 5.715 0.91 ;
        RECT 4.695 0.74 4.935 0.91 ;
        RECT 4.755 1.47 4.875 2.21 ;
        RECT 3.855 0.74 4.095 0.91 ;
        RECT 3.915 1.47 4.035 2.21 ;
        RECT 3.015 0.74 3.255 0.91 ;
        RECT 3.075 1.465 3.195 2.21 ;
        RECT 2.175 0.74 2.415 0.91 ;
        RECT 2.235 1.465 2.355 2.21 ;
        RECT 1.335 0.74 1.575 0.91 ;
        RECT 1.395 1.465 1.515 2.21 ;
        RECT 0.495 0.74 0.735 0.86 ;
        RECT 0.555 1.465 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 6.015 -0.18 6.135 0.67 ;
        RECT 5.175 -0.18 5.295 0.67 ;
        RECT 4.335 -0.18 4.455 0.67 ;
        RECT 3.495 -0.18 3.615 0.67 ;
        RECT 2.655 -0.18 2.775 0.67 ;
        RECT 1.815 -0.18 1.935 0.67 ;
        RECT 0.975 -0.18 1.095 0.665 ;
        RECT 0.135 -0.18 0.255 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 6.015 1.47 6.135 2.79 ;
        RECT 5.175 1.74 5.295 2.79 ;
        RECT 4.335 1.74 4.455 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
END INVX16

MACRO ADDHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX4 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 0.81 3.155 0.93 ;
        RECT 2.915 0.36 3.035 0.93 ;
        RECT 2.075 0.36 3.035 0.48 ;
        RECT 1.595 0.9 2.195 1.02 ;
        RECT 2.075 0.36 2.195 1.02 ;
        RECT 1.595 0.37 1.715 1.02 ;
        RECT 1.115 0.37 1.715 0.49 ;
        RECT 1.115 0.37 1.235 0.9 ;
        RECT 0.755 0.78 1.235 0.9 ;
        RECT 0.755 0.78 0.875 1.17 ;
        RECT 0.65 0.885 0.875 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.735 1.7 7.135 1.82 ;
        RECT 7.015 1.02 7.135 1.82 ;
        RECT 4.675 1.97 5.855 2.09 ;
        RECT 5.735 1.7 5.855 2.09 ;
        RECT 3.35 2.13 4.795 2.25 ;
        RECT 4.675 1.97 4.795 2.25 ;
        RECT 3.275 1.01 3.515 1.13 ;
        RECT 3.35 1.01 3.47 2.25 ;
        RECT 2.835 1.33 3.47 1.45 ;
        RECT 1.51 1.79 2.955 1.91 ;
        RECT 2.835 1.33 2.955 1.91 ;
        RECT 0.17 1.7 1.63 1.82 ;
        RECT 0.17 1.02 0.29 1.82 ;
        RECT 0.07 1.175 0.29 1.435 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.55 2.715 1.67 ;
        RECT 1.355 1.14 2.435 1.26 ;
        RECT 2.315 0.6 2.435 1.26 ;
        RECT 2.1 1.14 2.25 1.67 ;
        RECT 1.515 1.4 2.25 1.52 ;
        RECT 1.515 1.4 1.755 1.58 ;
        RECT 1.355 0.61 1.475 1.26 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.455 1.22 6.575 1.58 ;
        RECT 5.375 0.74 6.575 0.86 ;
        RECT 5.495 1.22 6.575 1.34 ;
        RECT 6.16 1.175 6.31 1.435 ;
        RECT 6.19 0.74 6.31 1.435 ;
        RECT 5.495 1.22 5.615 1.85 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 6.815 -0.18 7.055 0.38 ;
        RECT 5.915 -0.18 6.035 0.38 ;
        RECT 4.895 -0.18 5.135 0.38 ;
        RECT 3.155 -0.18 3.275 0.65 ;
        RECT 1.835 -0.18 1.955 0.78 ;
        RECT 0.875 -0.18 0.995 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.935 1.98 7.055 2.79 ;
        RECT 5.975 1.94 6.095 2.79 ;
        RECT 5.015 2.21 5.135 2.79 ;
        RECT 3.075 1.57 3.195 2.79 ;
        RECT 1.995 2.03 2.235 2.79 ;
        RECT 1.035 1.94 1.275 2.79 ;
        RECT 0.135 1.94 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.475 1.46 7.415 1.46 7.415 1.58 7.295 1.58 7.295 1.34 7.355 1.34 7.355 0.62 4.655 0.62 4.655 0.53 4.075 0.53 4.075 0.91 4.255 0.91 4.255 1.11 4.575 1.11 4.575 1.37 4.455 1.37 4.455 1.23 4.135 1.23 4.135 1.15 3.875 1.15 3.875 0.91 3.955 0.91 3.955 0.41 4.775 0.41 4.775 0.5 7.355 0.5 7.355 0.49 7.475 0.49 ;
      POLYGON 5.255 1.24 5.155 1.24 5.155 1.85 4.495 1.85 4.495 2.01 4.255 2.01 4.255 1.73 5.035 1.73 5.035 0.99 4.375 0.99 4.375 0.77 4.195 0.77 4.195 0.65 4.495 0.65 4.495 0.87 5.255 0.87 ;
      POLYGON 4.915 1.61 4.015 1.61 4.015 1.85 3.895 1.85 3.895 1.39 3.635 1.39 3.635 0.67 3.715 0.67 3.715 0.41 3.835 0.41 3.835 0.79 3.755 0.79 3.755 1.27 4.015 1.27 4.015 1.49 4.795 1.49 4.795 1.11 4.915 1.11 ;
      POLYGON 1.235 1.41 0.735 1.41 0.735 1.58 0.615 1.58 0.615 1.41 0.41 1.41 0.41 0.9 0.235 0.9 0.235 0.61 0.355 0.61 0.355 0.78 0.53 0.78 0.53 1.29 1.115 1.29 1.115 1.02 1.235 1.02 ;
  END
END ADDHX4

MACRO SDFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX8 0 0 ;
  SIZE 13.92 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.035 1.43 7.275 1.55 ;
        RECT 7.035 1.43 7.155 1.88 ;
        RECT 6.465 1.76 7.155 1.88 ;
        RECT 4.885 1.88 6.585 2 ;
        RECT 4.885 1.24 5.025 1.48 ;
        RECT 4.885 1.24 5.005 2 ;
        RECT 4.655 1.52 5.005 1.67 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.52 11.005 1.695 ;
        RECT 10.675 1.435 10.915 1.585 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.035 1.2 11.405 1.39 ;
        RECT 11.035 1.185 11.295 1.4 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.775 1.22 13.035 1.45 ;
        RECT 12.685 1.22 13.035 1.425 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.41 1.175 13.56 1.435 ;
        RECT 13.41 0.98 13.53 1.435 ;
        RECT 12.185 0.98 13.53 1.1 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5194 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 1.35 3.255 1.47 ;
        RECT 3.135 0.65 3.255 1.47 ;
        RECT 3.075 1.35 3.195 1.59 ;
        RECT 2.235 0.65 2.355 2.09 ;
        RECT 2.1 1.105 2.355 1.435 ;
        RECT 0.555 1.105 2.355 1.225 ;
        RECT 1.395 0.65 1.515 2.09 ;
        RECT 0.555 0.655 0.675 2.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.92 0.18 ;
        RECT 13.665 -0.18 13.785 0.4 ;
        RECT 12.805 -0.18 12.925 0.62 ;
        RECT 11.345 0.46 11.585 0.58 ;
        RECT 11.465 -0.18 11.585 0.58 ;
        RECT 10.145 0.465 10.385 0.585 ;
        RECT 10.265 -0.18 10.385 0.585 ;
        RECT 8.035 -0.18 8.155 0.73 ;
        RECT 6.855 -0.18 6.975 0.68 ;
        RECT 4.765 0.52 5.005 0.64 ;
        RECT 4.765 -0.18 4.885 0.64 ;
        RECT 3.985 -0.18 4.105 0.7 ;
        RECT 2.655 -0.18 2.775 0.64 ;
        RECT 1.815 -0.18 1.935 0.64 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.92 2.79 ;
        RECT 13.665 2.015 13.785 2.79 ;
        RECT 12.905 1.885 13.025 2.79 ;
        RECT 11.265 1.56 11.385 2.79 ;
        RECT 10.035 1.46 10.155 2.79 ;
        RECT 7.905 2.23 8.145 2.79 ;
        RECT 6.945 2.24 7.185 2.79 ;
        RECT 5.605 2.12 5.845 2.24 ;
        RECT 5.605 2.12 5.725 2.79 ;
        RECT 4.645 2.12 4.885 2.24 ;
        RECT 4.645 2.12 4.765 2.79 ;
        RECT 3.805 1.56 3.925 2.79 ;
        RECT 2.655 1.59 2.775 2.79 ;
        RECT 1.815 1.35 1.935 2.79 ;
        RECT 0.975 1.345 1.095 2.79 ;
        RECT 0.135 1.345 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.395 1.675 13.275 1.675 13.275 1.69 12.405 1.69 12.405 1.34 11.885 1.34 11.885 1.37 11.765 1.37 11.765 1.13 11.945 1.13 11.945 0.74 13.375 0.74 13.375 0.86 12.065 0.86 12.065 1.22 12.525 1.22 12.525 1.57 13.155 1.57 13.155 1.555 13.395 1.555 ;
      POLYGON 12.385 2.21 12.265 2.21 12.265 1.93 12.165 1.93 12.165 1.81 11.525 1.81 11.525 0.82 11.105 0.82 11.105 0.53 10.625 0.53 10.625 0.825 9.905 0.825 9.905 0.48 9.335 0.48 9.335 0.61 9.425 0.61 9.425 1.81 9.345 1.81 9.345 2.01 9.225 2.01 9.225 1.69 9.305 1.69 9.305 0.73 9.215 0.73 9.215 0.36 10.025 0.36 10.025 0.705 10.505 0.705 10.505 0.41 11.225 0.41 11.225 0.7 11.705 0.7 11.705 0.5 12.225 0.5 12.225 0.62 11.825 0.62 11.825 0.82 11.645 0.82 11.645 1.69 12.285 1.69 12.285 1.81 12.385 1.81 ;
      POLYGON 10.985 1.065 10.555 1.065 10.555 1.815 10.845 1.815 10.845 2.055 10.725 2.055 10.725 1.935 10.435 1.935 10.435 1.065 9.825 1.065 9.825 0.945 10.745 0.945 10.745 0.65 10.985 0.65 ;
      POLYGON 9.785 0.72 9.705 0.72 9.705 1.46 9.735 1.46 9.735 2.25 8.295 2.25 8.295 2.11 7.62 2.11 7.62 2.12 6.825 2.12 6.825 2.24 6.115 2.24 6.115 2.12 6.705 2.12 6.705 2 7.5 2 7.5 1.99 8.415 1.99 8.415 2.13 8.985 2.13 8.985 1.37 9.105 1.37 9.105 2.13 9.615 2.13 9.615 1.58 9.585 1.58 9.585 0.72 9.545 0.72 9.545 0.6 9.785 0.6 ;
      POLYGON 9.185 1.15 9.065 1.15 9.065 0.97 8.975 0.97 8.975 0.53 8.495 0.53 8.495 0.89 8.605 0.89 8.605 1.33 8.625 1.33 8.625 1.57 8.505 1.57 8.505 1.45 8.485 1.45 8.485 1.01 8.375 1.01 8.375 0.97 7.795 0.97 7.795 0.48 7.315 0.48 7.315 0.92 6.825 0.92 6.825 1.04 6.585 1.04 6.585 0.5 5.765 0.5 5.765 0.98 5.845 0.98 5.845 1.22 5.645 1.22 5.645 0.38 6.705 0.38 6.705 0.8 7.195 0.8 7.195 0.36 7.915 0.36 7.915 0.85 8.375 0.85 8.375 0.41 9.095 0.41 9.095 0.85 9.185 0.85 ;
      POLYGON 8.865 1.81 8.825 1.81 8.825 2.01 8.705 2.01 8.705 1.81 8.245 1.81 8.245 1.53 7.685 1.53 7.685 1.41 8.365 1.41 8.365 1.69 8.745 1.69 8.745 1.21 8.735 1.21 8.735 0.77 8.615 0.77 8.615 0.65 8.855 0.65 8.855 1.09 8.865 1.09 ;
      POLYGON 8.365 1.28 7.545 1.28 7.545 1.75 7.665 1.75 7.665 1.87 7.425 1.87 7.425 1.28 6.875 1.28 6.875 1.64 6.755 1.64 6.755 1.28 6.305 1.28 6.305 0.64 6.425 0.64 6.425 1.16 7.435 1.16 7.435 0.6 7.675 0.6 7.675 0.72 7.555 0.72 7.555 1.16 8.365 1.16 ;
      POLYGON 6.455 1.64 6.335 1.64 6.335 1.52 6.065 1.52 6.065 1.46 5.145 1.46 5.145 1.12 4.705 1.12 4.705 1.15 4.465 1.15 4.465 1 5.265 1 5.265 1.34 5.965 1.34 5.965 0.86 5.885 0.86 5.885 0.62 6.005 0.62 6.005 0.74 6.085 0.74 6.085 1.34 6.185 1.34 6.185 1.4 6.455 1.4 ;
      RECT 5.125 1.64 6.095 1.76 ;
      POLYGON 5.505 1.2 5.385 1.2 5.385 0.88 4.345 0.88 4.345 2.21 4.225 2.21 4.225 0.94 3.685 0.94 3.685 1.86 3.505 1.86 3.505 2.21 3.385 2.21 3.385 1.74 3.565 1.74 3.565 0.94 3.375 0.94 3.375 0.53 3.015 0.53 3.015 1.23 2.895 1.23 2.895 0.41 3.495 0.41 3.495 0.65 3.685 0.65 3.685 0.82 4.225 0.82 4.225 0.76 4.405 0.76 4.405 0.64 4.525 0.64 4.525 0.76 5.505 0.76 ;
  END
END SDFFSHQX8

MACRO DFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX2 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.115 0.9 7.235 1.31 ;
        RECT 6.975 0.9 7.235 1.13 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.165 1.475 1.38 ;
        RECT 1.185 1.14 1.47 1.38 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.23 3.175 1.38 ;
        RECT 2.595 1.36 3.035 1.48 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 1.465 0.8 1.725 ;
        RECT 0.645 1.4 0.77 1.725 ;
        RECT 0.645 0.68 0.765 2.05 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.385 -0.18 7.505 0.54 ;
        RECT 6.835 0.42 7.075 0.54 ;
        RECT 6.835 -0.18 6.955 0.54 ;
        RECT 4.975 0.43 5.215 0.55 ;
        RECT 5.095 -0.18 5.215 0.55 ;
        RECT 2.675 0.46 2.915 0.58 ;
        RECT 2.795 -0.18 2.915 0.58 ;
        RECT 1.005 0.66 1.245 0.78 ;
        RECT 1.005 -0.18 1.125 0.78 ;
        RECT 0.225 -0.18 0.345 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.445 2.23 7.565 2.79 ;
        RECT 5.655 2.26 5.895 2.79 ;
        RECT 4.575 2.01 4.815 2.13 ;
        RECT 4.575 2.01 4.695 2.79 ;
        RECT 2.975 1.84 3.095 2.79 ;
        RECT 2.855 1.84 3.095 1.96 ;
        RECT 1.875 1.74 1.995 2.79 ;
        RECT 1.065 1.5 1.185 2.79 ;
        RECT 0.225 1.4 0.345 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.985 1.81 7.865 1.81 7.865 1.55 6.825 1.55 6.825 1.43 7.355 1.43 7.355 0.78 6.56 0.78 6.56 0.48 6.015 0.48 6.015 0.92 6.135 0.92 6.135 1.04 5.895 1.04 5.895 0.79 4.735 0.79 4.735 0.48 4.095 0.48 4.095 0.92 4.375 0.92 4.375 1.04 3.975 1.04 3.975 0.36 4.855 0.36 4.855 0.67 5.895 0.67 5.895 0.36 6.68 0.36 6.68 0.66 7.475 0.66 7.475 1.43 7.865 1.43 7.865 0.4 7.985 0.4 ;
      POLYGON 7.905 2.25 7.785 2.25 7.785 2.11 7.11 2.11 7.11 2.25 6.195 2.25 6.195 2.14 4.935 2.14 4.935 1.89 3.975 1.89 3.975 2.23 3.295 2.23 3.295 1.72 2.735 1.72 2.735 2.25 2.115 2.25 2.115 1.62 1.605 1.62 1.605 1.74 1.485 1.74 1.485 1.5 1.605 1.5 1.605 0.6 1.725 0.6 1.725 1.5 2.235 1.5 2.235 2.13 2.615 2.13 2.615 1.6 3.295 1.6 3.295 1.06 3.175 1.06 3.175 0.94 3.415 0.94 3.415 2.11 3.855 2.11 3.855 1.33 3.775 1.33 3.775 1.21 4.015 1.21 4.015 1.33 3.975 1.33 3.975 1.77 5.055 1.77 5.055 2.02 6.345 2.02 6.345 1.52 6.225 1.52 6.225 1.4 6.465 1.4 6.465 2.13 6.99 2.13 6.99 1.99 7.905 1.99 ;
      POLYGON 6.705 2.01 6.585 2.01 6.585 1.28 4.855 1.28 4.855 1.39 4.735 1.39 4.735 1.15 4.855 1.15 4.855 1.16 6.255 1.16 6.255 0.72 6.135 0.72 6.135 0.6 6.375 0.6 6.375 1.16 6.705 1.16 ;
      POLYGON 6.225 1.9 6.105 1.9 6.105 1.87 5.415 1.87 5.415 1.9 5.175 1.9 5.175 1.75 6.105 1.75 6.105 1.66 6.225 1.66 ;
      POLYGON 5.775 1.04 5.535 1.04 5.535 1.03 4.615 1.03 4.615 1.65 4.095 1.65 4.095 1.53 4.495 1.53 4.495 0.72 4.215 0.72 4.215 0.6 4.615 0.6 4.615 0.91 5.655 0.91 5.655 0.92 5.775 0.92 ;
      POLYGON 3.735 1.99 3.615 1.99 3.615 1.59 3.535 1.59 3.535 0.82 2.455 0.82 2.455 1 2.175 1 2.175 0.88 2.335 0.88 2.335 0.7 3.535 0.7 3.535 0.5 3.655 0.5 3.655 1.47 3.735 1.47 ;
      POLYGON 3.055 1.11 2.695 1.11 2.695 1.24 2.475 1.24 2.475 2.01 2.355 2.01 2.355 1.24 1.935 1.24 1.935 0.6 2.095 0.6 2.095 0.48 1.485 0.48 1.485 1.02 1.025 1.02 1.025 1.26 0.905 1.26 0.905 0.9 1.365 0.9 1.365 0.36 2.215 0.36 2.215 0.72 2.055 0.72 2.055 1.12 2.575 1.12 2.575 0.99 3.055 0.99 ;
  END
END DFFRHQX2

MACRO DFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX4 0 0 ;
  SIZE 13.63 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.325 0.51 1.725 ;
        RECT 0.39 1.22 0.51 1.725 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 1.465 0.84 1.725 ;
        RECT 0.655 1.38 0.84 1.725 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 0.945 4.245 1.145 ;
        RECT 3.785 0.92 4.045 1.145 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 1.09 5.025 1.21 ;
        RECT 4.365 1.23 4.625 1.38 ;
        RECT 4.505 1.09 4.625 1.38 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.475 0.74 10.675 0.86 ;
        RECT 10.375 1.42 10.495 2.19 ;
        RECT 10.195 1.42 10.495 1.54 ;
        RECT 9.585 1.3 10.315 1.42 ;
        RECT 9.585 1.23 9.845 1.42 ;
        RECT 9.535 1.42 9.835 1.54 ;
        RECT 9.715 0.74 9.835 1.54 ;
        RECT 9.535 1.42 9.655 2.19 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.395 0.74 12.595 0.86 ;
        RECT 12.055 1.42 12.175 2.19 ;
        RECT 11.875 1.42 12.175 1.54 ;
        RECT 11.09 1.3 11.995 1.42 ;
        RECT 11.215 1.3 11.515 1.54 ;
        RECT 11.395 0.74 11.515 1.54 ;
        RECT 11.215 1.3 11.335 2.19 ;
        RECT 11.09 1.175 11.24 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.63 0.18 ;
        RECT 12.955 -0.18 13.075 0.73 ;
        RECT 11.875 -0.18 12.115 0.38 ;
        RECT 10.915 -0.18 11.155 0.38 ;
        RECT 9.955 -0.18 10.195 0.38 ;
        RECT 8.995 -0.18 9.115 0.82 ;
        RECT 8.155 -0.18 8.275 0.86 ;
        RECT 4.645 0.61 4.885 0.73 ;
        RECT 4.765 -0.18 4.885 0.73 ;
        RECT 2.095 -0.18 2.335 0.32 ;
        RECT 0.555 -0.18 0.675 0.86 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.63 2.79 ;
        RECT 12.475 1.54 12.595 2.79 ;
        RECT 11.635 1.54 11.755 2.79 ;
        RECT 10.795 1.54 10.915 2.79 ;
        RECT 9.955 1.54 10.075 2.79 ;
        RECT 9.115 1.64 9.235 2.79 ;
        RECT 8.275 1.7 8.395 2.79 ;
        RECT 7.155 1.88 7.395 2 ;
        RECT 7.155 1.88 7.275 2.79 ;
        RECT 3.985 2.22 4.225 2.79 ;
        RECT 2.805 2.225 3.045 2.79 ;
        RECT 1.895 2.225 2.015 2.79 ;
        RECT 0.555 1.92 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.495 0.92 13.335 0.92 13.335 1.42 13.015 1.42 13.015 2.19 12.895 2.19 12.895 1.42 12.295 1.42 12.295 1.28 12.535 1.28 12.535 1.3 13.215 1.3 13.215 0.8 13.375 0.8 13.375 0.68 13.495 0.68 ;
      POLYGON 13.095 1.18 12.855 1.18 12.855 0.97 12.715 0.97 12.715 0.62 9.355 0.62 9.355 1.06 8.855 1.06 8.855 1.18 9.455 1.18 9.455 1.3 8.855 1.3 8.855 1.76 8.815 1.76 8.815 2.16 8.695 2.16 8.695 1.64 8.735 1.64 8.735 1.22 7.615 1.22 7.615 1.1 8.575 1.1 8.575 0.68 8.695 0.68 8.695 0.94 9.235 0.94 9.235 0.5 12.835 0.5 12.835 0.85 12.975 0.85 12.975 1.06 13.095 1.06 ;
      POLYGON 8.615 1.52 6.265 1.52 6.265 1.71 6.025 1.71 6.025 0.67 6.145 0.67 6.145 1.4 8.375 1.4 8.375 1.36 8.615 1.36 ;
      POLYGON 8.035 1.88 7.515 1.88 7.515 1.76 6.445 1.76 6.445 1.64 7.635 1.64 7.635 1.76 8.035 1.76 ;
      POLYGON 7.855 0.86 7.735 0.86 7.735 0.56 7.075 0.56 7.075 0.8 6.835 0.8 6.835 0.68 6.955 0.68 6.955 0.44 7.855 0.44 ;
      POLYGON 7.495 0.8 7.315 0.8 7.315 1.04 6.595 1.04 6.595 0.91 6.505 0.91 6.505 0.67 6.625 0.67 6.625 0.79 6.715 0.79 6.715 0.92 7.195 0.92 7.195 0.68 7.495 0.68 ;
      POLYGON 7.235 1.28 6.355 1.28 6.355 1.15 6.265 1.15 6.265 0.55 5.305 0.55 5.305 1.53 5.065 1.53 5.065 1.41 5.185 1.41 5.185 0.97 4.39 0.97 4.39 0.48 4.085 0.48 4.085 0.36 4.51 0.36 4.51 0.85 5.185 0.85 5.185 0.43 6.385 0.43 6.385 1.03 6.475 1.03 6.475 1.16 7.235 1.16 ;
      POLYGON 7.025 2.05 6.785 2.05 6.785 2.01 4.585 2.01 4.585 1.86 3.765 1.86 3.765 1.625 2.765 1.625 2.765 1.22 2.885 1.22 2.885 1.505 3.885 1.505 3.885 1.74 4.705 1.74 4.705 1.89 5.785 1.89 5.785 1.17 5.665 1.17 5.665 1.05 5.905 1.05 5.905 1.89 6.905 1.89 6.905 1.93 7.025 1.93 ;
      POLYGON 6.005 2.25 4.345 2.25 4.345 2.1 3.525 2.1 3.525 1.865 2.435 1.865 2.435 1.745 2.525 1.745 2.525 1.46 1.535 1.46 1.535 1.32 1.775 1.32 1.775 1.34 2.525 1.34 2.525 0.72 2.765 0.72 2.765 0.84 2.645 0.84 2.645 1.745 3.645 1.745 3.645 1.98 4.465 1.98 4.465 2.13 6.005 2.13 ;
      POLYGON 5.725 0.93 5.545 0.93 5.545 1.53 5.665 1.53 5.665 1.77 4.825 1.77 4.825 1.62 4.005 1.62 4.005 1.385 3.545 1.385 3.545 1.1 2.885 1.1 2.885 0.56 1.855 0.56 1.855 0.48 1.735 0.48 1.735 0.36 1.975 0.36 1.975 0.44 3.005 0.44 3.005 0.98 3.545 0.98 3.545 0.8 3.485 0.8 3.485 0.68 3.725 0.68 3.725 0.8 3.665 0.8 3.665 1.265 4.245 1.265 4.245 1.5 4.945 1.5 4.945 1.65 5.425 1.65 5.425 0.81 5.605 0.81 5.605 0.67 5.725 0.67 ;
      POLYGON 4.165 0.8 3.845 0.8 3.845 0.56 3.365 0.56 3.365 0.62 3.245 0.62 3.245 0.86 3.125 0.86 3.125 0.5 3.245 0.5 3.245 0.44 3.965 0.44 3.965 0.68 4.165 0.68 ;
      POLYGON 3.405 2.25 3.165 2.25 3.165 2.105 1.195 2.105 1.195 1.84 1.295 1.84 1.295 0.96 1.255 0.96 1.255 0.62 1.375 0.62 1.375 0.84 1.415 0.84 1.415 1.985 3.285 1.985 3.285 2.13 3.405 2.13 ;
      POLYGON 2.405 1.22 2.285 1.22 2.285 1.06 1.695 1.06 1.695 1.18 1.575 1.18 1.575 0.72 1.495 0.72 1.495 0.5 1.135 0.5 1.135 1.48 1.175 1.48 1.175 1.72 1.015 1.72 1.015 1.1 0.24 1.1 0.24 1.845 0.255 1.845 0.255 2.085 0.135 2.085 0.135 1.965 0.12 1.965 0.12 0.86 0.135 0.86 0.135 0.62 0.255 0.62 0.255 0.98 1.015 0.98 1.015 0.38 1.615 0.38 1.615 0.6 1.695 0.6 1.695 0.94 2.405 0.94 ;
  END
END DFFNSRX4

MACRO TLATNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX4 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.14 0.52 1.59 ;
    END
  END GN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.19 0.4 4.755 0.52 ;
        RECT 2.13 0.5 3.31 0.62 ;
        RECT 2.13 0.36 2.25 0.62 ;
        RECT 1.355 0.36 2.25 0.48 ;
        RECT 0.655 1.16 1.475 1.28 ;
        RECT 1.355 0.36 1.475 1.28 ;
        RECT 1.175 1.16 1.435 1.38 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.465 2.67 1.585 ;
        RECT 2.55 1.335 2.67 1.585 ;
        RECT 2.39 1.465 2.54 1.73 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 1.15 6.395 1.27 ;
        RECT 5.815 1.15 6.075 1.38 ;
        RECT 5.255 1.36 5.935 1.48 ;
        RECT 5.255 1.17 5.375 1.48 ;
        RECT 5.095 1.17 5.375 1.29 ;
    END
  END SN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.855 1.31 7.975 2.08 ;
        RECT 7.675 1.31 7.975 1.43 ;
        RECT 7.035 0.85 7.815 0.97 ;
        RECT 7.695 0.68 7.815 0.97 ;
        RECT 7.03 1.19 7.795 1.31 ;
        RECT 7.03 1.175 7.18 1.435 ;
        RECT 7.035 0.8 7.155 1.435 ;
        RECT 7.015 1.31 7.135 2.08 ;
        RECT 6.855 0.8 7.155 0.92 ;
        RECT 6.855 0.68 6.975 0.92 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.215 1.31 11.335 2.08 ;
        RECT 11.035 1.31 11.335 1.43 ;
        RECT 10.395 0.85 11.175 0.97 ;
        RECT 11.055 0.68 11.175 0.97 ;
        RECT 10.395 1.19 11.155 1.31 ;
        RECT 10.395 0.85 10.715 1.31 ;
        RECT 10.375 1.31 10.515 1.43 ;
        RECT 10.375 1.31 10.495 2.08 ;
        RECT 10.215 0.8 10.515 0.92 ;
        RECT 10.215 0.68 10.335 0.92 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.475 -0.18 11.595 0.73 ;
        RECT 10.635 -0.18 10.755 0.73 ;
        RECT 9.795 -0.18 9.915 0.73 ;
        RECT 8.955 -0.18 9.075 0.73 ;
        RECT 8.115 -0.18 8.235 0.73 ;
        RECT 7.275 -0.18 7.395 0.73 ;
        RECT 6.435 -0.18 6.555 0.73 ;
        RECT 5.015 -0.18 5.135 0.8 ;
        RECT 2.915 -0.18 3.035 0.38 ;
        RECT 2.525 -0.18 2.645 0.38 ;
        RECT 0.555 -0.18 0.675 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 11.635 1.43 11.755 2.79 ;
        RECT 10.795 1.43 10.915 2.79 ;
        RECT 9.955 1.43 10.075 2.79 ;
        RECT 9.115 1.43 9.235 2.79 ;
        RECT 8.275 1.43 8.395 2.79 ;
        RECT 7.435 1.43 7.555 2.79 ;
        RECT 6.595 1.84 6.715 2.79 ;
        RECT 5.755 2.23 5.875 2.79 ;
        RECT 4.915 2.23 5.035 2.79 ;
        RECT 3.955 2 4.075 2.79 ;
        RECT 2.27 2.22 2.51 2.79 ;
        RECT 1.4 2.22 1.64 2.79 ;
        RECT 0.5 2.23 0.62 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.275 1.18 9.475 1.18 9.475 1.31 9.655 1.31 9.655 2.08 9.535 2.08 9.535 1.43 9.355 1.43 9.355 1.31 8.815 1.31 8.815 2.08 8.695 2.08 8.695 0.92 8.535 0.92 8.535 0.68 8.655 0.68 8.655 0.8 8.815 0.8 8.815 1.06 9.375 1.06 9.375 0.68 9.495 0.68 9.495 1.06 10.275 1.06 ;
      POLYGON 6.735 1.24 6.635 1.24 6.635 1.72 6.235 1.72 6.235 1.95 6.115 1.95 6.115 1.72 5.395 1.72 5.395 1.95 5.275 1.95 5.275 1.72 4.855 1.72 4.855 1.45 4.295 1.45 4.295 1.33 4.975 1.33 4.975 1.6 6.515 1.6 6.515 1.03 5.735 1.03 5.735 0.66 5.855 0.66 5.855 0.91 6.735 0.91 ;
      POLYGON 5.615 1.24 5.495 1.24 5.495 1.04 4.175 1.04 4.175 1.64 3.23 1.64 3.23 1.82 3.15 1.82 3.15 1.94 3.03 1.94 3.03 1.7 3.11 1.7 3.11 1.52 4.055 1.52 4.055 1.04 3.695 1.04 3.695 0.92 3.615 0.92 3.615 0.66 3.735 0.66 3.735 0.8 3.815 0.8 3.815 0.92 5.615 0.92 ;
      RECT 3.39 1.76 4.615 1.88 ;
      POLYGON 3.935 1.28 3.815 1.28 3.815 1.4 2.99 1.4 2.99 1.58 2.91 1.58 2.91 1.97 2.27 1.97 2.27 2.1 1.55 2.1 1.55 1.62 1.1 1.62 1.1 1.83 0.98 1.83 0.98 1.5 1.595 1.5 1.595 0.6 1.835 0.6 1.835 0.72 1.715 0.72 1.715 1.62 1.67 1.62 1.67 1.98 2.15 1.98 2.15 1.225 2.39 1.225 2.39 1.345 2.27 1.345 2.27 1.85 2.79 1.85 2.79 1.28 3.695 1.28 3.695 1.16 3.935 1.16 ;
      POLYGON 3.575 1.16 3.335 1.16 3.335 1.105 2.03 1.105 2.03 1.86 1.79 1.86 1.79 1.74 1.91 1.74 1.91 0.84 1.985 0.84 1.985 0.74 2.225 0.74 2.225 0.985 3.455 0.985 3.455 1.04 3.575 1.04 ;
      POLYGON 1.235 1.04 0.995 1.04 0.995 1.02 0.24 1.02 0.24 1.71 0.255 1.71 0.255 1.95 0.135 1.95 0.135 1.83 0.12 1.83 0.12 0.78 0.135 0.78 0.135 0.54 0.255 0.54 0.255 0.9 1.235 0.9 ;
  END
END TLATNSRX4

MACRO ADDFHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX2 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.505 0.83 6.545 0.95 ;
        RECT 4.565 0.82 4.685 1.06 ;
        RECT 3.205 0.78 3.625 0.9 ;
        RECT 3.205 0.65 3.465 0.9 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.325 1.07 7.445 1.31 ;
        RECT 5.095 1.07 7.445 1.19 ;
        RECT 6.975 0.94 7.235 1.19 ;
        RECT 4.325 1.18 5.215 1.3 ;
        RECT 3.065 1.07 4.445 1.19 ;
        RECT 2.8 1.02 3.185 1.14 ;
        RECT 2.005 0.99 2.92 1.11 ;
        RECT 1.885 1.06 2.125 1.18 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.335 1.31 7.165 1.43 ;
        RECT 2.915 1.42 5.455 1.54 ;
        RECT 2.915 1.31 3.175 1.67 ;
        RECT 2.79 1.31 3.175 1.43 ;
        RECT 2.285 1.26 2.91 1.35 ;
        RECT 2.525 1.31 3.175 1.38 ;
        RECT 2.285 1.23 2.645 1.35 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.585 0.68 0.705 2.21 ;
        RECT 0.36 0.885 0.705 1.145 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.025 0.885 8.34 1.145 ;
        RECT 8.025 0.59 8.145 1.68 ;
        RECT 7.905 1.56 8.025 2.21 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 8.445 -0.18 8.565 0.64 ;
        RECT 7.485 0.35 7.725 0.47 ;
        RECT 7.485 -0.18 7.605 0.47 ;
        RECT 5.065 0.35 5.305 0.47 ;
        RECT 5.065 -0.18 5.185 0.47 ;
        RECT 4.225 -0.18 4.345 0.64 ;
        RECT 1.965 -0.18 2.205 0.38 ;
        RECT 1.005 -0.18 1.125 0.73 ;
        RECT 0.165 -0.18 0.285 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 8.325 1.56 8.445 2.79 ;
        RECT 7.425 2.03 7.665 2.15 ;
        RECT 7.425 2.03 7.545 2.79 ;
        RECT 5.225 2.23 5.345 2.79 ;
        RECT 4.205 2.22 4.445 2.79 ;
        RECT 1.965 2.2 2.205 2.79 ;
        RECT 1.065 1.98 1.185 2.79 ;
        RECT 0.165 1.56 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.885 1.44 7.685 1.44 7.685 1.91 6.605 1.91 6.605 2.21 6.485 2.21 6.485 1.91 6.185 1.91 6.185 2.07 6.065 2.07 6.065 1.79 7.565 1.79 7.565 0.71 6.085 0.71 6.085 0.63 5.965 0.63 5.965 0.51 6.205 0.51 6.205 0.59 6.625 0.59 6.625 0.45 6.745 0.45 6.745 0.59 7.685 0.59 7.685 1.2 7.885 1.2 ;
      POLYGON 6.425 1.67 5.945 1.67 5.945 2.11 4.89 2.11 4.89 2.1 3.685 2.1 3.685 2.2 3.565 2.2 3.565 2.1 2.925 2.1 2.925 2.08 1.51 2.08 1.51 1.86 1.245 1.86 1.245 1.26 0.825 1.26 0.825 1.14 1.245 1.14 1.245 0.5 2.925 0.5 2.925 0.41 3.585 0.41 3.585 0.4 3.705 0.4 3.705 0.64 3.585 0.64 3.585 0.53 3.045 0.53 3.045 0.82 2.925 0.82 2.925 0.62 1.365 0.62 1.365 1.74 1.63 1.74 1.63 1.96 2.925 1.96 2.925 1.79 3.045 1.79 3.045 1.98 3.565 1.98 3.565 1.68 3.685 1.68 3.685 1.98 5.01 1.98 5.01 1.99 5.825 1.99 5.825 1.55 6.425 1.55 ;
      POLYGON 5.725 0.71 4.805 0.71 4.805 0.68 4.585 0.68 4.585 0.56 4.925 0.56 4.925 0.59 5.605 0.59 5.605 0.47 5.725 0.47 ;
      POLYGON 5.705 1.87 5.585 1.87 5.585 1.86 4.685 1.86 4.685 1.74 5.585 1.74 5.585 1.55 5.705 1.55 ;
      RECT 1.485 0.74 2.685 0.86 ;
      POLYGON 2.685 1.84 2.445 1.84 2.445 1.62 1.665 1.62 1.665 1.34 1.785 1.34 1.785 1.5 2.565 1.5 2.565 1.57 2.685 1.57 ;
  END
END ADDFHX2

MACRO OR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.395 1.32 ;
        RECT 0.275 1.08 0.395 1.32 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.39 1.09 1.725 ;
        RECT 0.815 1.39 1.09 1.625 ;
        RECT 0.815 1.29 0.935 1.625 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.485 0.68 1.605 0.92 ;
        RECT 1.395 0.8 1.515 1.965 ;
        RECT 1.23 1.465 1.515 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 1.035 -0.18 1.155 0.4 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.845 1.095 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.255 1.27 1.135 1.27 1.135 1.17 0.675 1.17 0.675 1.905 0.275 1.905 0.275 1.785 0.555 1.785 0.555 0.68 0.675 0.68 0.675 1.05 1.135 1.05 1.135 1.03 1.255 1.03 ;
  END
END OR2XL

MACRO NOR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X6 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.415 0.99 4.535 1.26 ;
        RECT 0.68 0.99 4.535 1.11 ;
        RECT 3.175 0.99 3.415 1.195 ;
        RECT 1.955 0.99 2.195 1.195 ;
        RECT 0.65 1.08 0.8 1.435 ;
        RECT 0.435 1.08 0.8 1.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.3 4.235 1.42 ;
        RECT 3.785 1.23 4.045 1.42 ;
        RECT 1.315 1.315 3.905 1.435 ;
        RECT 2.315 1.3 2.555 1.435 ;
        RECT 1.195 1.3 1.435 1.42 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.4496 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.555 4.775 1.675 ;
        RECT 4.655 0.75 4.775 1.675 ;
        RECT 4.42 1.465 4.775 1.675 ;
        RECT 0.555 0.75 4.775 0.87 ;
        RECT 4.42 1.465 4.57 1.725 ;
        RECT 3.935 1.555 4.055 2.21 ;
        RECT 3.915 0.4 4.035 0.87 ;
        RECT 3.075 0.4 3.195 0.87 ;
        RECT 2.495 1.555 2.615 2.21 ;
        RECT 2.235 0.4 2.355 0.87 ;
        RECT 1.395 0.4 1.515 0.87 ;
        RECT 1.175 1.555 1.295 2.21 ;
        RECT 0.555 0.4 0.675 0.87 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.275 0.46 4.515 0.63 ;
        RECT 4.275 -0.18 4.395 0.63 ;
        RECT 3.435 0.46 3.675 0.63 ;
        RECT 3.435 -0.18 3.555 0.63 ;
        RECT 2.595 0.46 2.835 0.63 ;
        RECT 2.595 -0.18 2.715 0.63 ;
        RECT 1.755 0.46 1.995 0.63 ;
        RECT 1.755 -0.18 1.875 0.63 ;
        RECT 0.915 0.46 1.155 0.63 ;
        RECT 0.915 -0.18 1.035 0.63 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 4.575 1.845 4.695 2.79 ;
        RECT 3.295 1.795 3.415 2.79 ;
        RECT 1.815 1.795 1.935 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
END NOR2X6

MACRO NOR2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.24 3.615 1.48 ;
        RECT 3.29 1.36 3.615 1.48 ;
        RECT 3.26 1.465 3.41 1.725 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.25 2.555 1.37 ;
        RECT 2.045 1.23 2.305 1.38 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9664 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.73 3.195 0.85 ;
        RECT 3.075 0.61 3.195 0.85 ;
        RECT 2.355 1.5 2.475 2.21 ;
        RECT 2.235 0.61 2.355 0.85 ;
        RECT 0.175 1.5 2.475 1.62 ;
        RECT 1.395 0.61 1.515 0.85 ;
        RECT 1.075 1.5 1.195 2.21 ;
        RECT 0.555 0.61 0.675 0.85 ;
        RECT 0.175 1.23 0.565 1.38 ;
        RECT 0.175 0.73 0.295 1.62 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.495 -0.18 3.615 0.85 ;
        RECT 2.595 0.48 2.835 0.6 ;
        RECT 2.595 -0.18 2.715 0.6 ;
        RECT 1.755 0.48 1.995 0.6 ;
        RECT 1.755 -0.18 1.875 0.6 ;
        RECT 0.915 0.48 1.155 0.6 ;
        RECT 0.915 -0.18 1.035 0.6 ;
        RECT 0.075 0.48 0.315 0.6 ;
        RECT 0.075 -0.18 0.195 0.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.295 1.845 3.415 2.79 ;
        RECT 1.715 1.74 1.835 2.79 ;
        RECT 0.335 1.74 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.035 0.99 3.895 0.99 3.895 1.8 3.775 1.8 3.775 1.11 3.335 1.11 3.335 1.13 3.095 1.13 3.095 1.11 1.925 1.11 1.925 1.13 1.685 1.13 1.685 1.11 0.415 1.11 0.415 0.99 3.775 0.99 3.775 0.87 3.915 0.87 3.915 0.61 4.035 0.61 ;
  END
END NOR2BX4

MACRO AOI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 0.82 1.96 1.16 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 1.315 1.38 1.725 ;
        RECT 1.21 1.3 1.33 1.725 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.465 1.01 1.625 ;
        RECT 0.89 1.385 1.01 1.625 ;
        RECT 0.65 1.465 0.8 1.725 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.52 0.81 0.64 ;
        RECT 0.25 0.82 0.69 0.94 ;
        RECT 0.57 0.52 0.69 0.94 ;
        RECT 0.41 1.3 0.53 1.965 ;
        RECT 0.07 1.3 0.53 1.42 ;
        RECT 0.07 1.175 0.37 1.42 ;
        RECT 0.25 0.82 0.37 1.42 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.89 -0.18 2.01 0.7 ;
        RECT 1.05 -0.18 1.17 0.7 ;
        RECT 0.21 -0.18 0.33 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.05 1.845 1.17 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.87 1.905 1.5 1.905 1.5 1.18 0.49 1.18 0.49 1.06 1.5 1.06 1.5 0.7 1.47 0.7 1.47 0.46 1.59 0.46 1.59 0.58 1.62 0.58 1.62 1.785 1.87 1.785 ;
  END
END AOI2BB1XL

MACRO NOR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X8 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.695 0.81 9.815 1.21 ;
        RECT 9.005 0.81 9.815 0.93 ;
        RECT 1.855 0.73 9.125 0.845 ;
        RECT 6.035 0.81 9.815 0.85 ;
        RECT 7.15 1.03 7.39 1.15 ;
        RECT 7.15 0.73 7.27 1.15 ;
        RECT 1.855 0.725 6.155 0.845 ;
        RECT 4.465 1.03 4.705 1.15 ;
        RECT 4.585 0.725 4.705 1.15 ;
        RECT 1.855 0.725 2.015 1.09 ;
        RECT 1.735 1.035 1.975 1.155 ;
        RECT 1.755 0.94 2.015 1.09 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.23 9.555 1.38 ;
        RECT 9.295 1.05 9.535 1.38 ;
        RECT 8.765 1.05 9.535 1.17 ;
        RECT 7.97 0.97 8.885 1.09 ;
        RECT 7.65 1.05 8.155 1.17 ;
        RECT 6.855 1.27 7.77 1.39 ;
        RECT 7.65 1.05 7.77 1.39 ;
        RECT 6.855 1.05 6.975 1.39 ;
        RECT 5.795 1.05 6.975 1.17 ;
        RECT 5.195 0.965 5.915 1.085 ;
        RECT 4.825 1.05 5.315 1.17 ;
        RECT 4.225 1.27 4.945 1.39 ;
        RECT 4.825 1.05 4.945 1.39 ;
        RECT 4.225 0.99 4.345 1.39 ;
        RECT 3.695 0.99 4.345 1.11 ;
        RECT 3.695 0.965 3.815 1.23 ;
        RECT 2.9 0.965 3.815 1.085 ;
        RECT 2.135 1.055 3.02 1.175 ;
        RECT 1.405 1.275 2.255 1.395 ;
        RECT 2.135 1.055 2.255 1.395 ;
        RECT 1.405 1.055 1.525 1.395 ;
        RECT 0.755 1.055 1.525 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 1.21 8.555 1.33 ;
        RECT 8.315 1.21 8.435 1.63 ;
        RECT 2.565 1.51 8.435 1.63 ;
        RECT 5.435 1.205 5.675 1.325 ;
        RECT 5.435 1.205 5.555 1.63 ;
        RECT 3.355 1.205 3.475 1.63 ;
        RECT 3.235 1.205 3.475 1.325 ;
        RECT 0.975 1.515 2.685 1.635 ;
        RECT 0.975 1.295 1.095 1.635 ;
        RECT 0.445 1.295 1.095 1.415 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.445 1.125 0.565 1.415 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.6308 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.495 0.485 10.335 0.605 ;
        RECT 9.835 1.52 10.135 1.67 ;
        RECT 1.835 1.755 10.055 1.875 ;
        RECT 9.935 0.485 10.055 1.875 ;
        RECT 9.835 1.47 9.955 2.21 ;
        RECT 7.49 1.75 7.61 2.21 ;
        RECT 4.245 1.75 4.365 2.21 ;
        RECT 1.835 1.755 1.955 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 9.615 -0.18 9.855 0.365 ;
        RECT 8.655 -0.18 8.895 0.365 ;
        RECT 7.695 -0.18 7.935 0.365 ;
        RECT 6.735 -0.18 6.975 0.365 ;
        RECT 5.775 -0.18 6.015 0.365 ;
        RECT 4.815 -0.18 5.055 0.365 ;
        RECT 3.855 -0.18 4.095 0.365 ;
        RECT 2.895 -0.18 3.135 0.365 ;
        RECT 1.935 -0.18 2.175 0.365 ;
        RECT 0.975 -0.18 1.215 0.365 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 8.595 1.995 8.835 2.15 ;
        RECT 8.595 1.995 8.715 2.79 ;
        RECT 5.515 1.995 5.755 2.15 ;
        RECT 5.515 1.995 5.635 2.79 ;
        RECT 2.955 1.995 3.195 2.15 ;
        RECT 2.955 1.995 3.075 2.79 ;
        RECT 0.335 1.535 0.455 2.79 ;
    END
  END VDD
END NOR3X8

MACRO ADDHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX2 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.075 0.42 5.315 0.54 ;
        RECT 3.485 0.5 5.195 0.62 ;
        RECT 1.255 0.48 3.605 0.6 ;
        RECT 3.215 0.38 3.455 0.6 ;
        RECT 2.815 0.48 2.935 1.46 ;
        RECT 0.535 0.645 1.375 0.765 ;
        RECT 1.255 0.48 1.375 0.765 ;
        RECT 0.535 0.885 0.8 1.145 ;
        RECT 0.535 0.645 0.655 1.24 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.54 1.94 2.66 2.24 ;
        RECT 2.38 1.94 2.66 2.06 ;
        RECT 1.315 1.86 2.5 1.98 ;
        RECT 1.315 1.3 1.435 1.98 ;
        RECT 1.175 1.3 1.435 1.67 ;
        RECT 1.16 1.3 1.435 1.42 ;
    END
  END A
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 1.465 1.96 1.725 ;
        RECT 1.66 1.62 1.92 1.74 ;
        RECT 1.8 0.72 1.92 1.74 ;
        RECT 1.495 0.72 1.92 0.84 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.355 0.885 4.57 1.145 ;
        RECT 4.32 1.4 4.56 1.52 ;
        RECT 4.355 0.74 4.475 1.52 ;
        RECT 4.235 0.74 4.475 0.86 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.715 -0.18 4.955 0.38 ;
        RECT 3.755 -0.18 3.995 0.38 ;
        RECT 1.975 -0.18 2.215 0.36 ;
        RECT 1.015 -0.18 1.135 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.8 2.04 5.04 2.16 ;
        RECT 4.8 2.04 4.92 2.79 ;
        RECT 3.84 1.88 4.08 2 ;
        RECT 3.84 1.88 3.96 2.79 ;
        RECT 2.2 2.22 2.32 2.79 ;
        RECT 1.18 2.1 1.42 2.22 ;
        RECT 1.18 2.1 1.3 2.79 ;
        RECT 0.34 1.68 0.46 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.435 0.86 5.375 0.86 5.375 1.76 3.93 1.76 3.93 1.48 3.295 1.48 3.295 1.24 3.415 1.24 3.415 1.36 4.05 1.36 4.05 1.64 5.255 1.64 5.255 0.86 5.195 0.86 5.195 0.74 5.435 0.74 ;
      POLYGON 4.22 1.24 4.1 1.24 4.1 1.12 3.175 1.12 3.175 1.7 3.16 1.7 3.16 1.82 3.04 1.82 3.04 1.58 3.055 1.58 3.055 0.72 3.295 0.72 3.295 0.84 3.175 0.84 3.175 1 4.22 1 ;
      POLYGON 3.72 2.18 2.78 2.18 2.78 1.82 2.62 1.82 2.62 1.7 2.575 1.7 2.575 0.84 2.455 0.84 2.455 0.72 2.695 0.72 2.695 1.58 2.74 1.58 2.74 1.7 2.9 1.7 2.9 2.06 3.72 2.06 ;
      POLYGON 1.68 1.3 1.56 1.3 1.56 1.18 1.04 1.18 1.04 1.74 0.7 1.74 0.7 1.62 0.92 1.62 0.92 1.48 0.295 1.48 0.295 0.66 0.415 0.66 0.415 1.36 0.92 1.36 0.92 1.06 1.68 1.06 ;
  END
END ADDHX2

MACRO OR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X6 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.06 1.635 1.18 ;
        RECT 0.36 1.175 0.56 1.3 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.3 1.015 1.42 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.3 0.8 1.725 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.235 0.91 4.095 1.03 ;
        RECT 3.975 0.4 4.095 1.03 ;
        RECT 3.775 1.39 3.895 2.21 ;
        RECT 2.095 1.39 3.895 1.51 ;
        RECT 3.175 0.885 3.41 1.145 ;
        RECT 3.175 0.795 3.295 1.51 ;
        RECT 3.135 0.4 3.255 1.03 ;
        RECT 2.935 1.39 3.055 2.21 ;
        RECT 2.235 0.4 2.355 1.03 ;
        RECT 2.095 1.39 2.215 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.555 -0.18 3.675 0.79 ;
        RECT 2.715 -0.18 2.835 0.79 ;
        RECT 1.815 -0.18 1.935 0.7 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.355 1.63 3.475 2.79 ;
        RECT 2.515 1.63 2.635 2.79 ;
        RECT 1.675 1.56 1.795 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.055 1.27 1.875 1.27 1.875 1.44 1.255 1.44 1.255 1.68 1.095 1.68 1.095 2.21 0.975 2.21 0.975 1.56 1.135 1.56 1.135 1.32 1.755 1.32 1.755 0.94 0.555 0.94 0.555 0.59 0.675 0.59 0.675 0.82 1.395 0.82 1.395 0.59 1.515 0.59 1.515 0.82 1.875 0.82 1.875 1.15 3.055 1.15 ;
  END
END OR2X6

MACRO OAI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.06 3.315 1.18 ;
        RECT 2.39 1.06 2.54 1.435 ;
        RECT 2.115 1.18 2.54 1.3 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.97 1.755 1.21 ;
        RECT 1.465 0.94 1.725 1.09 ;
        RECT 0.415 0.97 1.755 1.09 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.465 3.12 1.725 ;
        RECT 2.97 1.3 3.09 1.725 ;
        RECT 2.735 1.3 3.09 1.42 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.28 1.155 1.4 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.28 0.8 1.725 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.015 0.65 3.255 0.77 ;
        RECT 2.15 0.76 3.135 0.88 ;
        RECT 2.655 1.555 2.775 2.21 ;
        RECT 1.135 1.555 2.775 1.675 ;
        RECT 2.15 0.65 2.415 0.88 ;
        RECT 1.875 0.94 2.27 1.06 ;
        RECT 2.15 0.65 2.27 1.06 ;
        RECT 1.755 1.52 2.015 1.675 ;
        RECT 1.875 0.94 1.995 1.675 ;
        RECT 1.135 1.555 1.255 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 1.335 0.46 1.575 0.58 ;
        RECT 1.335 -0.18 1.455 0.58 ;
        RECT 0.495 0.46 0.735 0.58 ;
        RECT 0.495 -0.18 0.615 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.295 1.56 3.415 2.79 ;
        RECT 1.855 1.795 2.095 2.15 ;
        RECT 1.855 1.795 1.975 2.79 ;
        RECT 0.495 1.845 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.615 0.65 3.495 0.65 3.495 0.53 2.775 0.53 2.775 0.64 2.655 0.64 2.655 0.53 1.935 0.53 1.935 0.82 0.195 0.82 0.195 0.77 0.075 0.77 0.075 0.65 0.315 0.65 0.315 0.7 0.915 0.7 0.915 0.65 1.155 0.65 1.155 0.7 1.815 0.7 1.815 0.41 2.655 0.41 2.655 0.4 2.775 0.4 2.775 0.41 3.615 0.41 ;
  END
END OAI22X2

MACRO CLKBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX8 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.87 0.825 3.99 1.305 ;
        RECT 3.84 0.825 3.99 1.28 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.69 0.715 2.93 0.835 ;
        RECT 2.75 1.295 2.87 2.21 ;
        RECT 0.23 0.76 2.81 0.88 ;
        RECT 2.57 1.295 2.87 1.415 ;
        RECT 0.23 1.27 2.69 1.39 ;
        RECT 1.85 0.71 2.09 0.88 ;
        RECT 1.91 1.27 2.03 2.21 ;
        RECT 1.01 0.71 1.25 0.88 ;
        RECT 1.07 1.27 1.19 2.21 ;
        RECT 0.36 0.76 0.51 1.145 ;
        RECT 0.36 0.76 0.48 1.39 ;
        RECT 0.23 1.27 0.35 2.21 ;
        RECT 0.23 0.64 0.35 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 4.01 -0.18 4.13 0.705 ;
        RECT 3.17 -0.18 3.29 0.705 ;
        RECT 2.33 -0.18 2.45 0.64 ;
        RECT 1.49 -0.18 1.61 0.64 ;
        RECT 0.65 -0.18 0.77 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 4.01 1.465 4.13 2.79 ;
        RECT 3.17 1.465 3.29 2.79 ;
        RECT 2.33 1.51 2.45 2.79 ;
        RECT 1.49 1.51 1.61 2.79 ;
        RECT 0.65 1.51 0.77 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.71 2.115 3.59 2.115 3.59 1.15 3.19 1.15 3.19 1.175 2.95 1.175 2.95 1.15 0.87 1.15 0.87 1.03 3.59 1.03 3.59 0.655 3.71 0.655 ;
  END
END CLKBUFX8

MACRO TLATNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX1 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.845 1.3 2.165 1.42 ;
        RECT 1.81 1.465 1.965 1.725 ;
        RECT 1.845 1.3 1.965 1.725 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.175 5.15 1.51 ;
        RECT 4.915 1.24 5.035 1.57 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.67 1.4 6.91 1.52 ;
        RECT 6.245 1.36 6.79 1.48 ;
        RECT 6.105 1.23 6.375 1.38 ;
        RECT 6.255 0.48 6.375 1.48 ;
        RECT 5.265 0.48 6.375 0.6 ;
        RECT 4.725 0.5 5.385 0.62 ;
        RECT 3.015 0.4 4.845 0.52 ;
    END
  END RN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.155 1.28 7.275 1.565 ;
        RECT 7.03 1.43 7.18 1.725 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 2.21 ;
        RECT 1.23 1.175 1.485 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 6.995 -0.18 7.115 0.92 ;
        RECT 5.025 -0.18 5.145 0.38 ;
        RECT 2.775 0.72 3.115 0.84 ;
        RECT 2.775 -0.18 2.895 0.84 ;
        RECT 1.785 -0.18 1.905 0.73 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.995 1.845 7.115 2.79 ;
        RECT 6.155 1.845 6.275 2.79 ;
        RECT 5.075 1.7 5.195 2.79 ;
        RECT 3.585 2.07 3.705 2.79 ;
        RECT 2.745 2.23 2.865 2.79 ;
        RECT 1.785 1.845 1.905 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.535 1.965 7.415 1.965 7.415 1.16 6.615 1.16 6.615 1.24 6.495 1.24 6.495 1 6.615 1 6.615 1.04 7.415 1.04 7.415 0.68 7.535 0.68 ;
      POLYGON 6.695 1.965 6.575 1.965 6.575 1.845 6.43 1.845 6.43 1.725 5.865 1.725 5.865 1.34 5.51 1.34 5.51 1.22 5.865 1.22 5.865 0.74 6.135 0.74 6.135 0.86 5.985 0.86 5.985 1.605 6.55 1.605 6.55 1.725 6.695 1.725 ;
      POLYGON 5.745 0.84 5.625 0.84 5.625 1.055 5.39 1.055 5.39 1.46 5.615 1.46 5.615 1.82 5.495 1.82 5.495 1.58 5.27 1.58 5.27 1.055 4.795 1.055 4.795 1.38 3.975 1.38 3.975 1.26 4.595 1.26 4.595 1.02 4.675 1.02 4.675 0.935 5.505 0.935 5.505 0.72 5.745 0.72 ;
      POLYGON 4.555 0.9 4.475 0.9 4.475 1.14 3.855 1.14 3.855 1.5 4.435 1.5 4.435 1.82 4.315 1.82 4.315 1.62 3.735 1.62 3.735 1.51 2.545 1.51 2.545 1.27 2.665 1.27 2.665 1.39 3.735 1.39 3.735 1.02 4.355 1.02 4.355 0.78 4.435 0.78 4.435 0.66 4.555 0.66 ;
      RECT 3.045 1.74 4.075 1.86 ;
      POLYGON 3.615 1.16 3.375 1.16 3.375 1.15 2.405 1.15 2.405 1.66 2.385 1.66 2.385 1.83 2.265 1.83 2.265 1.54 2.285 1.54 2.285 1.15 1.725 1.15 1.725 1.27 1.605 1.27 1.605 1.03 2.485 1.03 2.485 0.68 2.605 0.68 2.605 1.03 3.615 1.03 ;
      POLYGON 1.095 1.99 0.975 1.99 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END TLATNSRX1

MACRO NAND4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BXL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.85 0.51 1.35 ;
        RECT 0.36 0.85 0.51 1.32 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.905 0.935 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.885 1.38 1.275 ;
        RECT 1.14 0.83 1.26 1.23 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.72 1.175 2.015 1.445 ;
        RECT 1.72 1.175 1.96 1.46 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2976 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 1.65 1.575 1.77 ;
        RECT 1.335 1.47 1.455 1.77 ;
        RECT 0.12 1.47 1.455 1.59 ;
        RECT 0.495 1.47 0.735 1.77 ;
        RECT 0.07 0.595 0.455 0.73 ;
        RECT 0.335 0.49 0.455 0.73 ;
        RECT 0.12 0.595 0.24 1.59 ;
        RECT 0.07 0.595 0.24 0.855 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.62 -0.18 1.74 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.875 2.23 1.995 2.79 ;
        RECT 0.915 2.23 1.035 2.79 ;
        RECT 0.135 1.71 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.475 1.83 2.355 1.83 2.355 1.71 2.135 1.71 2.135 1.01 1.5 1.01 1.5 0.89 2.135 0.89 2.135 0.73 2.04 0.73 2.04 0.49 2.16 0.49 2.16 0.61 2.255 0.61 2.255 1.59 2.475 1.59 ;
  END
END NAND4BXL

MACRO TLATNCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX16 0 0 ;
  SIZE 13.92 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.845 0.8 1.145 ;
        RECT 0.555 0.975 0.675 1.26 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.83 1.175 13.1 1.435 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.335 0.74 6.575 0.86 ;
        RECT 5.555 0.79 6.455 0.91 ;
        RECT 6.075 1.49 6.315 1.61 ;
        RECT 1.295 1.37 6.195 1.49 ;
        RECT 5.555 0.67 5.675 1.49 ;
        RECT 5.235 1.37 5.475 1.61 ;
        RECT 4.655 0.74 4.895 0.86 ;
        RECT 4.71 1.175 4.86 1.49 ;
        RECT 4.395 1.37 4.83 1.61 ;
        RECT 4.71 0.74 4.83 1.61 ;
        RECT 3.695 0.74 4.055 0.86 ;
        RECT 3.495 1.37 3.815 1.61 ;
        RECT 3.695 0.74 3.815 1.61 ;
        RECT 2.795 0.74 3.215 0.86 ;
        RECT 2.655 1.37 2.915 1.61 ;
        RECT 2.795 0.74 2.915 1.61 ;
        RECT 1.955 0.74 2.315 0.86 ;
        RECT 1.815 1.37 2.075 1.61 ;
        RECT 1.955 0.74 2.075 1.61 ;
        RECT 0.975 1.49 1.415 1.61 ;
        RECT 1.295 0.68 1.415 1.61 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.92 0.18 ;
        RECT 13.07 0.455 13.31 0.575 ;
        RECT 13.19 -0.18 13.31 0.575 ;
        RECT 11.095 -0.18 11.215 0.49 ;
        RECT 10.135 -0.18 10.255 0.67 ;
        RECT 8.415 0.37 8.655 0.49 ;
        RECT 8.415 -0.18 8.535 0.49 ;
        RECT 6.815 -0.18 6.935 0.67 ;
        RECT 5.975 -0.18 6.095 0.67 ;
        RECT 5.135 -0.18 5.255 0.67 ;
        RECT 4.295 -0.18 4.415 0.67 ;
        RECT 3.455 -0.18 3.575 0.67 ;
        RECT 2.555 -0.18 2.675 0.665 ;
        RECT 1.715 -0.18 1.835 0.665 ;
        RECT 0.875 -0.18 0.995 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.92 2.79 ;
        RECT 13.07 1.635 13.19 2.79 ;
        RECT 11.23 2.055 11.47 2.175 ;
        RECT 11.23 2.055 11.35 2.79 ;
        RECT 10.395 2.23 10.515 2.79 ;
        RECT 9.375 1.97 9.615 2.09 ;
        RECT 9.375 1.97 9.495 2.79 ;
        RECT 8.415 1.97 8.655 2.09 ;
        RECT 8.415 1.97 8.535 2.79 ;
        RECT 7.455 1.97 7.695 2.09 ;
        RECT 7.455 1.97 7.575 2.79 ;
        RECT 6.495 1.97 6.735 2.11 ;
        RECT 6.495 1.97 6.615 2.79 ;
        RECT 5.655 1.97 5.895 2.11 ;
        RECT 5.655 1.97 5.775 2.79 ;
        RECT 4.815 1.97 5.055 2.11 ;
        RECT 4.815 1.97 4.935 2.79 ;
        RECT 3.915 1.97 4.155 2.115 ;
        RECT 3.915 1.97 4.035 2.79 ;
        RECT 3.075 1.97 3.315 2.115 ;
        RECT 3.075 1.97 3.195 2.79 ;
        RECT 2.235 1.97 2.475 2.115 ;
        RECT 2.235 1.97 2.355 2.79 ;
        RECT 1.395 1.97 1.635 2.115 ;
        RECT 1.395 1.97 1.515 2.79 ;
        RECT 0.555 1.97 0.795 2.115 ;
        RECT 0.555 1.97 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.73 1.635 13.61 1.635 13.61 1.755 13.49 1.755 13.49 1.515 13.61 1.515 13.61 0.815 12.83 0.815 12.83 0.5 11.77 0.5 11.77 0.73 10.855 0.73 10.855 0.5 10.495 0.5 10.495 0.97 9.275 0.97 9.275 1.12 9.035 1.12 9.035 0.97 8.035 0.97 8.035 1.12 7.795 1.12 7.795 0.85 10.375 0.85 10.375 0.38 10.975 0.38 10.975 0.61 11.65 0.61 11.65 0.38 12.01 0.38 12.01 0.36 12.25 0.36 12.25 0.38 12.95 0.38 12.95 0.695 13.61 0.695 13.61 0.62 13.73 0.62 ;
      POLYGON 13.35 1.2 13.23 1.2 13.23 1.055 12.71 1.055 12.71 1.935 9.94 1.935 9.94 1.85 0.135 1.85 0.135 1.43 0.315 1.43 0.315 0.68 0.435 0.68 0.435 1.55 0.255 1.55 0.255 1.73 10.06 1.73 10.06 1.815 12.59 1.815 12.59 1.415 11.87 1.415 11.87 1.175 11.99 1.175 11.99 1.295 12.59 1.295 12.59 0.935 13.35 0.935 ;
      POLYGON 12.47 0.97 11.75 0.97 11.75 1.535 12.05 1.535 12.05 1.575 12.17 1.575 12.17 1.695 11.93 1.695 11.93 1.655 11.63 1.655 11.63 1.42 11.05 1.42 11.05 1.09 11.17 1.09 11.17 1.3 11.63 1.3 11.63 0.85 12.35 0.85 12.35 0.62 12.47 0.62 ;
      POLYGON 11.51 1.18 11.39 1.18 11.39 0.97 10.735 0.97 10.735 1.36 10.93 1.36 10.93 1.695 10.81 1.695 10.81 1.48 10.615 1.48 10.615 1.36 6.955 1.36 6.955 1.11 7.075 1.11 7.075 1.24 8.255 1.24 8.255 1.09 8.375 1.09 8.375 1.24 10.115 1.24 10.115 1.11 10.235 1.11 10.235 1.24 10.615 1.24 10.615 0.62 10.735 0.62 10.735 0.85 11.51 0.85 ;
      POLYGON 10.095 1.61 9.855 1.61 9.855 1.6 9.135 1.6 9.135 1.61 8.895 1.61 8.895 1.6 8.175 1.6 8.175 1.61 7.935 1.61 7.935 1.6 7.215 1.6 7.215 1.61 6.975 1.61 6.975 1.6 6.715 1.6 6.715 1.18 6.195 1.18 6.195 1.06 6.715 1.06 6.715 0.86 7.46 0.86 7.46 0.61 9.555 0.61 9.555 0.73 7.58 0.73 7.58 0.98 6.835 0.98 6.835 1.48 9.975 1.48 9.975 1.49 10.095 1.49 ;
  END
END TLATNCAX16

MACRO FILL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL1 0 0 ;
  SIZE 0.29 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.29 0.18 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.29 2.79 ;
    END
  END VDD
END FILL1

MACRO DFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX2 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.98 0.88 5.1 1.24 ;
        RECT 4.61 0.88 5.1 1 ;
        RECT 4.61 0.36 4.73 1 ;
        RECT 2.68 0.36 4.73 0.48 ;
        RECT 2.68 0.885 2.83 1.145 ;
        RECT 2.68 0.36 2.8 1.34 ;
        RECT 2.26 1.22 2.8 1.34 ;
        RECT 2.14 1.26 2.38 1.38 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.12 7.525 1.39 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.165 8.105 1.39 ;
        RECT 7.72 1.165 8.105 1.365 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.64 0.8 1.99 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.52 -0.18 7.64 0.74 ;
        RECT 5.88 -0.18 6.12 0.32 ;
        RECT 4.85 0.64 5.09 0.76 ;
        RECT 4.85 -0.18 4.97 0.76 ;
        RECT 1.94 -0.18 2.06 0.68 ;
        RECT 1.1 -0.18 1.22 0.69 ;
        RECT 0.26 -0.18 0.38 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.4 1.75 7.52 2.79 ;
        RECT 6.06 1.68 6.18 2.79 ;
        RECT 5.94 1.68 6.18 1.93 ;
        RECT 4.92 2.29 5.16 2.79 ;
        RECT 2.72 1.98 2.96 2.15 ;
        RECT 2.72 1.98 2.84 2.79 ;
        RECT 1.94 1.74 2.06 2.79 ;
        RECT 1.1 1.34 1.22 2.79 ;
        RECT 0.26 1.34 0.38 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.06 1 7.145 1 7.145 1.51 7.81 1.51 7.81 1.66 7.94 1.66 7.94 1.9 7.82 1.9 7.82 1.78 7.69 1.78 7.69 1.63 7.28 1.63 7.28 2.23 6.68 2.23 6.68 2.25 6.44 2.25 6.44 2.13 6.48 2.13 6.48 1.56 5.82 1.56 5.82 2.17 4.6 2.17 4.6 2.05 5.7 2.05 5.7 1.44 6.6 1.44 6.6 2.11 7.025 2.11 7.025 1 6.96 1 6.96 0.88 7.94 0.88 7.94 0.5 8.06 0.5 ;
      POLYGON 6.86 0.76 6.84 0.76 6.84 1.99 6.72 1.99 6.72 1.32 5.7 1.32 5.7 1.2 6.72 1.2 6.72 0.64 6.74 0.64 6.74 0.5 6.86 0.5 ;
      POLYGON 6.6 1.08 6.48 1.08 6.48 0.84 6.215 0.84 6.215 0.56 5.34 0.56 5.34 1.48 4.66 1.48 4.66 1.69 4.37 1.69 4.37 1.14 4.23 1.14 4.23 0.9 4.37 0.9 4.37 0.76 4.25 0.76 4.25 0.64 4.49 0.64 4.49 1.36 5.22 1.36 5.22 0.44 6.335 0.44 6.335 0.72 6.6 0.72 ;
      POLYGON 6.34 1.08 5.58 1.08 5.58 1.93 4.21 1.93 4.21 2.21 4.09 2.21 4.09 1.38 3.99 1.38 3.99 0.72 3.61 0.72 3.61 0.6 4.11 0.6 4.11 1.26 4.21 1.26 4.21 1.81 5.46 1.81 5.46 0.96 5.55 0.96 5.55 0.68 5.67 0.68 5.67 0.96 6.34 0.96 ;
      POLYGON 3.87 1.36 3.75 1.36 3.75 1.24 3.19 1.24 3.19 0.88 3.31 0.88 3.31 1.12 3.87 1.12 ;
      POLYGON 3.79 2.21 3.67 2.21 3.67 1.6 3.07 1.6 3.07 1.62 1.8 1.62 1.8 1.37 1.92 1.37 1.92 1.5 2.95 1.5 2.95 0.64 3.19 0.64 3.19 0.6 3.43 0.6 3.43 0.72 3.31 0.72 3.31 0.76 3.07 0.76 3.07 1.48 3.79 1.48 ;
      POLYGON 3.37 2.21 3.25 2.21 3.25 1.86 2.48 1.86 2.48 2.21 2.36 2.21 2.36 1.74 3.25 1.74 3.25 1.72 3.37 1.72 ;
      POLYGON 2.56 1.1 1.64 1.1 1.64 2.21 1.52 2.21 1.52 1.1 1.06 1.1 1.06 1.22 0.94 1.22 0.94 0.98 1.52 0.98 1.52 0.54 1.64 0.54 1.64 0.98 2.44 0.98 2.44 0.86 2.56 0.86 ;
  END
END DFFSHQX2

MACRO TBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX3 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 1.29 1.12 ;
        RECT 0.39 0.885 0.51 1.24 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.845 0.96 3 1.2 ;
        RECT 2.88 0.44 3 1.2 ;
        RECT 1.41 0.44 3 0.56 ;
        RECT 1.465 1.23 1.725 1.38 ;
        RECT 1.41 0.44 1.53 1.36 ;
        RECT 0.71 1.24 1.725 1.36 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.385 1.56 4.505 2.21 ;
        RECT 4.38 0.62 4.5 0.86 ;
        RECT 3.84 1.56 4.505 1.68 ;
        RECT 4.2 0.74 4.5 0.86 ;
        RECT 3.84 0.86 4.32 0.98 ;
        RECT 3.84 1.465 3.99 1.725 ;
        RECT 3.425 1.8 3.96 1.92 ;
        RECT 3.84 0.79 3.96 1.92 ;
        RECT 3.54 0.79 3.96 0.91 ;
        RECT 3.54 0.62 3.66 0.91 ;
        RECT 3.425 1.8 3.545 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.96 -0.18 4.08 0.67 ;
        RECT 3.12 -0.18 3.24 0.67 ;
        RECT 2.04 -0.18 2.28 0.32 ;
        RECT 0.93 -0.18 1.05 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.905 2.04 4.025 2.79 ;
        RECT 3.005 1.8 3.125 2.79 ;
        RECT 0.975 2.1 1.215 2.22 ;
        RECT 0.975 2.1 1.095 2.79 ;
        RECT 0.135 1.72 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.72 1.68 2.885 1.68 2.885 1.8 2.725 1.8 2.725 2.25 2.075 2.25 2.075 1.98 0.675 1.98 0.675 2.21 0.555 2.21 0.555 1.6 0.12 1.6 0.12 0.645 0.29 0.645 0.29 0.525 0.41 0.525 0.41 0.765 0.24 0.765 0.24 1.48 0.675 1.48 0.675 1.86 2.195 1.86 2.195 2.13 2.605 2.13 2.605 1.68 2.765 1.68 2.765 1.56 3.6 1.56 3.6 1.22 3.72 1.22 ;
      POLYGON 3.38 1.44 2.645 1.44 2.645 1.56 2.485 1.56 2.485 2.01 2.365 2.01 2.365 1.44 2.525 1.44 2.525 0.8 2.52 0.8 2.52 0.68 2.76 0.68 2.76 0.8 2.645 0.8 2.645 1.32 3.26 1.32 3.26 0.94 3.38 0.94 ;
      POLYGON 2.405 1.32 1.965 1.32 1.965 1.62 1.695 1.62 1.695 1.74 1.455 1.74 1.455 1.62 1.575 1.62 1.575 1.5 1.845 1.5 1.845 0.8 1.65 0.8 1.65 0.68 1.965 0.68 1.965 1.2 2.405 1.2 ;
  END
END TBUFX3

MACRO NOR2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX2 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.465 1.38 1.725 ;
        RECT 1.23 1.34 1.35 1.725 ;
        RECT 1.215 1.22 1.335 1.46 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1.24 2.015 1.585 ;
        RECT 1.81 1.465 1.96 1.725 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.69 1.575 0.81 ;
        RECT 0.175 0.74 1.455 0.86 ;
        RECT 0.975 1.32 1.095 2.21 ;
        RECT 0.175 1.32 1.095 1.44 ;
        RECT 0.495 0.69 0.735 0.86 ;
        RECT 0.07 1.175 0.295 1.435 ;
        RECT 0.175 0.74 0.295 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.815 -0.18 1.935 0.86 ;
        RECT 0.915 0.5 1.155 0.62 ;
        RECT 0.915 -0.18 1.035 0.62 ;
        RECT 0.075 0.5 0.315 0.62 ;
        RECT 0.075 -0.18 0.195 0.62 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.695 1.845 1.815 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.355 0.98 2.295 0.98 2.295 1.8 2.175 1.8 2.175 1.1 1.715 1.1 1.715 1.15 1.475 1.15 1.475 1.1 0.655 1.1 0.655 1.13 0.415 1.13 0.415 1.01 0.535 1.01 0.535 0.98 2.175 0.98 2.175 0.86 2.235 0.86 2.235 0.62 2.355 0.62 ;
  END
END NOR2BX2

MACRO AOI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X4 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.015 0.99 4.755 1.11 ;
        RECT 4.075 0.94 4.335 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.175 3.41 1.435 ;
        RECT 3.255 0.99 3.38 1.18 ;
        RECT 3.255 0.94 3.375 1.18 ;
        RECT 0.915 0.99 3.38 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.23 2.775 1.35 ;
        RECT 1.175 1.23 1.435 1.38 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9664 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.835 1.315 4.955 2.01 ;
        RECT 4.595 0.65 4.835 0.77 ;
        RECT 3.775 1.315 4.955 1.435 ;
        RECT 1.535 0.7 4.715 0.82 ;
        RECT 3.995 1.315 4.115 2.01 ;
        RECT 3.775 1.23 4.045 1.435 ;
        RECT 3.815 0.58 3.935 0.82 ;
        RECT 3.775 0.7 3.895 1.435 ;
        RECT 2.695 0.65 2.935 0.82 ;
        RECT 1.415 0.65 1.655 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 5.075 -0.18 5.195 0.64 ;
        RECT 4.175 0.46 4.415 0.58 ;
        RECT 4.175 -0.18 4.295 0.58 ;
        RECT 3.335 0.46 3.575 0.58 ;
        RECT 3.335 -0.18 3.455 0.58 ;
        RECT 2.055 0.46 2.295 0.58 ;
        RECT 2.055 -0.18 2.175 0.58 ;
        RECT 0.835 -0.18 0.955 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 3.095 1.795 3.335 2.15 ;
        RECT 3.095 1.795 3.215 2.79 ;
        RECT 2.255 1.795 2.495 2.15 ;
        RECT 2.255 1.795 2.375 2.79 ;
        RECT 1.415 1.795 1.655 2.15 ;
        RECT 1.415 1.795 1.535 2.79 ;
        RECT 0.575 1.795 0.815 2.15 ;
        RECT 0.575 1.795 0.695 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.375 2.25 3.575 2.25 3.575 1.675 2.855 1.675 2.855 2.21 2.735 2.21 2.735 1.675 2.015 1.675 2.015 2.21 1.895 2.21 1.895 1.675 1.175 1.675 1.175 2.21 1.055 2.21 1.055 1.675 0.335 1.675 0.335 2.21 0.215 2.21 0.215 1.555 3.695 1.555 3.695 2.13 4.415 2.13 4.415 1.56 4.535 1.56 4.535 2.13 5.255 2.13 5.255 1.56 5.375 1.56 ;
  END
END AOI21X4

MACRO SDFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX2 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.085 1.43 4.325 1.55 ;
        RECT 3.175 1.76 4.205 1.88 ;
        RECT 4.085 1.43 4.205 1.88 ;
        RECT 3.175 1.76 3.295 2.01 ;
        RECT 2.835 1.89 3.295 2.01 ;
        RECT 1.825 1.99 2.955 2.11 ;
        RECT 1.775 1.23 2.015 1.47 ;
        RECT 1.825 1.23 1.945 2.11 ;
        RECT 1.755 1.23 2.015 1.38 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.405 8.155 1.65 ;
        RECT 7.845 1.405 8.105 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 1.055 8.515 1.265 ;
        RECT 8.135 0.94 8.395 1.175 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.855 1.22 10.135 1.415 ;
        RECT 9.855 1.22 9.975 1.555 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 0.885 10.66 1.145 ;
        RECT 10.51 0.885 10.63 1.165 ;
        RECT 9.235 0.98 10.66 1.1 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.68 0.675 1.99 ;
        RECT 0.305 0.94 0.675 1.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.745 -0.18 10.865 0.765 ;
        RECT 9.855 -0.18 9.975 0.62 ;
        RECT 8.375 0.46 8.615 0.58 ;
        RECT 8.495 -0.18 8.615 0.58 ;
        RECT 7.175 -0.18 7.415 0.38 ;
        RECT 5.185 -0.18 5.305 0.75 ;
        RECT 4.005 -0.18 4.125 0.68 ;
        RECT 1.755 0.51 1.995 0.63 ;
        RECT 1.755 -0.18 1.875 0.63 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.745 1.475 10.865 2.79 ;
        RECT 10.015 1.915 10.135 2.79 ;
        RECT 8.515 1.56 8.635 2.79 ;
        RECT 7.175 1.46 7.295 2.79 ;
        RECT 4.865 2.23 5.105 2.79 ;
        RECT 3.905 2.24 4.145 2.79 ;
        RECT 2.545 2.23 2.785 2.79 ;
        RECT 1.585 2.23 1.825 2.79 ;
        RECT 0.975 1.34 1.095 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.505 0.705 10.385 0.705 10.385 0.86 9.115 0.86 9.115 1.3 9.735 1.3 9.735 1.675 10.265 1.675 10.265 1.535 10.505 1.535 10.505 1.655 10.385 1.655 10.385 1.795 9.615 1.795 9.615 1.42 8.995 1.42 8.995 1.09 8.875 1.09 8.875 0.97 8.995 0.97 8.995 0.74 10.265 0.74 10.265 0.585 10.505 0.585 ;
      POLYGON 9.495 2.21 9.375 2.21 9.375 1.66 8.755 1.66 8.755 1.44 8.635 1.44 8.635 0.82 8.135 0.82 8.135 0.53 7.655 0.53 7.655 0.62 6.485 0.62 6.485 1.75 6.505 1.75 6.505 2.01 6.265 2.01 6.265 1.75 6.365 1.75 6.365 0.5 7.535 0.5 7.535 0.41 8.255 0.41 8.255 0.7 8.75 0.7 8.75 0.5 9.255 0.5 9.255 0.62 8.87 0.62 8.87 0.82 8.755 0.82 8.755 1.32 8.875 1.32 8.875 1.54 9.495 1.54 ;
      POLYGON 8.015 0.86 7.725 0.86 7.725 1.79 7.955 1.79 7.955 2.03 7.835 2.03 7.835 1.91 7.605 1.91 7.605 1.19 6.975 1.19 6.975 1.07 7.605 1.07 7.605 0.74 7.775 0.74 7.775 0.65 8.015 0.65 ;
      POLYGON 6.935 0.86 6.855 0.86 6.855 1.46 6.875 1.46 6.875 2.25 5.495 2.25 5.495 2.11 4.595 2.11 4.595 2.12 3.535 2.12 3.535 2.25 3.075 2.25 3.075 2.13 3.415 2.13 3.415 2 4.475 2 4.475 1.99 5.615 1.99 5.615 2.13 6.025 2.13 6.025 1.37 6.145 1.37 6.145 2.13 6.755 2.13 6.755 1.58 6.735 1.58 6.735 0.86 6.695 0.86 6.695 0.74 6.935 0.74 ;
      POLYGON 6.245 1.17 6.125 1.17 6.125 0.55 5.645 0.55 5.645 1.27 5.665 1.27 5.665 1.39 5.425 1.39 5.425 1.27 5.525 1.27 5.525 0.99 4.945 0.99 4.945 0.48 4.465 0.48 4.465 0.92 3.895 0.92 3.895 1.04 3.655 1.04 3.655 0.92 3.695 0.92 3.695 0.48 2.755 0.48 2.755 0.96 2.835 0.96 2.835 1.2 2.635 1.2 2.635 0.36 3.815 0.36 3.815 0.8 4.345 0.8 4.345 0.36 5.065 0.36 5.065 0.87 5.525 0.87 5.525 0.43 6.245 0.43 ;
      POLYGON 6.005 0.79 5.905 0.79 5.905 1.63 5.855 1.63 5.855 2.01 5.735 2.01 5.735 1.63 4.705 1.63 4.705 1.35 4.825 1.35 4.825 1.51 5.785 1.51 5.785 0.79 5.765 0.79 5.765 0.67 6.005 0.67 ;
      POLYGON 5.305 1.23 4.565 1.23 4.565 1.75 4.625 1.75 4.625 1.87 4.385 1.87 4.385 1.75 4.445 1.75 4.445 1.23 4.135 1.23 4.135 1.31 3.835 1.31 3.835 1.64 3.715 1.64 3.715 1.28 3.415 1.28 3.415 0.84 3.295 0.84 3.295 0.6 3.415 0.6 3.415 0.72 3.535 0.72 3.535 1.16 4.015 1.16 4.015 1.11 4.585 1.11 4.585 0.6 4.825 0.6 4.825 0.72 4.705 0.72 4.705 1.11 5.305 1.11 ;
      POLYGON 3.415 1.64 3.295 1.64 3.295 1.52 3.175 1.52 3.175 1.44 2.135 1.44 2.135 1.11 1.455 1.11 1.455 0.99 2.255 0.99 2.255 1.32 2.955 1.32 2.955 0.84 2.875 0.84 2.875 0.6 2.995 0.6 2.995 0.72 3.075 0.72 3.075 1.32 3.295 1.32 3.295 1.4 3.415 1.4 ;
      POLYGON 3.055 1.77 2.305 1.77 2.305 1.87 2.065 1.87 2.065 1.75 2.185 1.75 2.185 1.65 2.815 1.65 2.815 1.56 3.055 1.56 ;
      POLYGON 2.495 1.16 2.375 1.16 2.375 0.87 1.335 0.87 1.335 1.34 1.515 1.34 1.515 1.86 1.395 1.86 1.395 1.46 1.215 1.46 1.215 1.2 0.795 1.2 0.795 1.08 1.215 1.08 1.215 0.71 1.395 0.71 1.395 0.59 1.515 0.59 1.515 0.75 2.495 0.75 ;
  END
END SDFFSHQX2

MACRO OAI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X4 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.155 0.82 4.275 1.15 ;
        RECT 2.31 0.82 4.275 0.94 ;
        RECT 1.895 0.97 2.43 1.09 ;
        RECT 2.045 0.94 2.43 1.09 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.14 8.215 1.38 ;
        RECT 6.755 1.06 8.055 1.18 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.35 1.27 5.315 1.39 ;
        RECT 3.35 1.06 3.47 1.39 ;
        RECT 2.555 1.06 3.47 1.18 ;
        RECT 1.015 1.21 2.675 1.33 ;
        RECT 2.555 1.06 2.675 1.33 ;
        RECT 1.175 1.21 1.435 1.38 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 1.175 8.63 1.435 ;
        RECT 6.175 1.5 8.6 1.62 ;
        RECT 8.435 1.24 8.6 1.62 ;
        RECT 7.375 1.3 7.615 1.62 ;
        RECT 6.175 1.22 6.295 1.62 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 1.51 5.655 1.63 ;
        RECT 5.535 1.24 5.655 1.63 ;
        RECT 2.99 1.3 3.23 1.63 ;
        RECT 0.735 1.23 0.855 1.63 ;
        RECT 0.595 1.23 0.855 1.38 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.815 0.65 9.055 0.77 ;
        RECT 6.295 0.76 8.935 0.88 ;
        RECT 7.975 0.65 8.215 0.88 ;
        RECT 7.935 1.74 8.055 2.21 ;
        RECT 1.875 1.75 8.055 1.87 ;
        RECT 7.135 0.65 7.375 0.88 ;
        RECT 6.655 1.74 6.775 2.21 ;
        RECT 6.295 0.65 6.535 0.88 ;
        RECT 5.935 0.82 6.415 0.94 ;
        RECT 5.815 1.75 6.075 1.96 ;
        RECT 5.935 0.82 6.055 1.96 ;
        RECT 4.435 1.75 4.555 2.21 ;
        RECT 1.875 1.75 1.995 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 5.395 0.34 5.635 0.46 ;
        RECT 5.395 -0.18 5.515 0.46 ;
        RECT 4.435 0.34 4.675 0.46 ;
        RECT 4.435 -0.18 4.555 0.46 ;
        RECT 3.475 0.34 3.715 0.46 ;
        RECT 3.475 -0.18 3.595 0.46 ;
        RECT 2.515 0.34 2.755 0.46 ;
        RECT 2.515 -0.18 2.635 0.46 ;
        RECT 1.555 0.34 1.795 0.46 ;
        RECT 1.555 -0.18 1.675 0.46 ;
        RECT 0.595 0.34 0.835 0.46 ;
        RECT 0.595 -0.18 0.715 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.575 1.74 8.695 2.79 ;
        RECT 7.235 1.99 7.475 2.15 ;
        RECT 7.235 1.99 7.355 2.79 ;
        RECT 5.815 2.08 6.055 2.2 ;
        RECT 5.815 2.08 5.935 2.79 ;
        RECT 3.27 1.99 3.51 2.15 ;
        RECT 3.27 1.99 3.39 2.79 ;
        RECT 0.595 1.75 0.715 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.415 0.65 9.295 0.65 9.295 0.53 8.575 0.53 8.575 0.64 8.455 0.64 8.455 0.53 7.735 0.53 7.735 0.64 7.615 0.64 7.615 0.53 6.895 0.53 6.895 0.64 6.775 0.64 6.775 0.53 6.055 0.53 6.055 0.7 0.115 0.7 0.115 0.58 5.935 0.58 5.935 0.41 6.775 0.41 6.775 0.4 6.895 0.4 6.895 0.41 7.615 0.41 7.615 0.4 7.735 0.4 7.735 0.41 8.455 0.41 8.455 0.4 8.575 0.4 8.575 0.41 9.415 0.41 ;
  END
END OAI32X4

MACRO CLKBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX12 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.45 1.3 4.775 1.42 ;
        RECT 4.42 1.465 4.57 1.725 ;
        RECT 4.45 1.3 4.57 1.725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.915 1.32 4.035 2.21 ;
        RECT 0.515 0.82 4.035 0.94 ;
        RECT 3.915 0.4 4.035 0.94 ;
        RECT 0.515 1.32 4.035 1.44 ;
        RECT 3.075 1.32 3.195 2.21 ;
        RECT 3.075 0.4 3.195 0.94 ;
        RECT 2.235 1.32 2.355 2.21 ;
        RECT 2.235 0.4 2.355 0.94 ;
        RECT 1.395 1.32 1.515 2.21 ;
        RECT 1.395 0.4 1.515 0.94 ;
        RECT 0.555 1.32 0.8 1.725 ;
        RECT 0.555 1.32 0.675 2.21 ;
        RECT 0.555 0.4 0.675 0.94 ;
        RECT 0.515 0.8 0.635 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.175 -0.18 5.295 0.725 ;
        RECT 4.335 -0.18 4.455 0.915 ;
        RECT 3.495 -0.18 3.615 0.7 ;
        RECT 2.655 -0.18 2.775 0.7 ;
        RECT 1.815 -0.18 1.935 0.7 ;
        RECT 0.975 -0.18 1.095 0.7 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.175 1.56 5.295 2.79 ;
        RECT 4.335 1.845 4.455 2.79 ;
        RECT 3.495 1.56 3.615 2.79 ;
        RECT 2.655 1.56 2.775 2.79 ;
        RECT 1.815 1.56 1.935 2.79 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.43 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.715 0.965 5.015 0.965 5.015 1.32 5.715 1.32 5.715 2.21 5.595 2.21 5.595 1.44 5.015 1.44 5.015 1.66 4.875 1.66 4.875 2.21 4.755 2.21 4.755 1.54 4.895 1.54 4.895 1.18 3.935 1.18 3.935 1.195 3.695 1.195 3.695 1.18 3.095 1.18 3.095 1.195 2.855 1.195 2.855 1.18 2.675 1.18 2.675 1.195 2.435 1.195 2.435 1.18 1.835 1.18 1.835 1.195 1.595 1.195 1.595 1.18 0.995 1.18 0.995 1.2 0.755 1.2 0.755 1.08 0.875 1.08 0.875 1.06 4.755 1.06 4.755 0.675 4.875 0.675 4.875 0.845 5.595 0.845 5.595 0.675 5.715 0.675 ;
  END
END CLKBUFX12

MACRO SDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX4 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.2 1.21 1.44 ;
        RECT 0.36 1.2 1.21 1.32 ;
        RECT 0.36 1.175 0.51 1.435 ;
        RECT 0.39 1.08 0.51 1.435 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 1.44 0.89 1.76 ;
        RECT 0.65 1.465 0.8 1.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.99 1.96 1.45 ;
        RECT 1.84 0.965 1.96 1.45 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.455 2.595 1.67 ;
        RECT 2.215 1.455 2.595 1.645 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.025 0.7 9.225 0.82 ;
        RECT 9.085 1.44 9.205 2.21 ;
        RECT 8.905 1.44 9.205 1.56 ;
        RECT 8.22 1.32 9.025 1.44 ;
        RECT 8.245 0.7 8.365 2.21 ;
        RECT 8.19 1.175 8.365 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.945 0.7 11.145 0.82 ;
        RECT 10.765 1.32 10.885 2.21 ;
        RECT 9.93 1.32 10.885 1.44 ;
        RECT 9.96 0.7 10.08 1.56 ;
        RECT 9.925 1.44 10.045 2.21 ;
        RECT 9.93 1.175 10.08 1.56 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.505 -0.18 11.625 0.69 ;
        RECT 10.425 -0.18 10.665 0.34 ;
        RECT 9.465 -0.18 9.705 0.34 ;
        RECT 8.505 -0.18 8.745 0.34 ;
        RECT 7.545 -0.18 7.785 0.34 ;
        RECT 6.705 -0.18 6.825 0.86 ;
        RECT 4.985 0.55 5.225 0.67 ;
        RECT 4.985 -0.18 5.105 0.67 ;
        RECT 2.935 -0.18 3.055 0.92 ;
        RECT 1.95 -0.18 2.07 0.845 ;
        RECT 0.615 -0.18 0.735 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.185 1.56 11.305 2.79 ;
        RECT 10.345 1.56 10.465 2.79 ;
        RECT 9.505 1.56 9.625 2.79 ;
        RECT 8.665 1.56 8.785 2.79 ;
        RECT 7.825 1.56 7.945 2.79 ;
        RECT 6.925 1.58 7.045 2.79 ;
        RECT 5.225 1.75 5.345 2.79 ;
        RECT 3.33 2.29 3.57 2.79 ;
        RECT 2.13 2.05 2.37 2.17 ;
        RECT 2.13 2.05 2.25 2.79 ;
        RECT 0.71 1.95 0.83 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.045 0.88 11.865 0.88 11.865 1.44 11.725 1.44 11.725 2.21 11.605 2.21 11.605 1.44 11.005 1.44 11.005 1.3 11.245 1.3 11.245 1.32 11.745 1.32 11.745 0.76 11.925 0.76 11.925 0.64 12.045 0.64 ;
      POLYGON 11.585 1.2 11.465 1.2 11.465 0.93 11.265 0.93 11.265 0.58 7.245 0.58 7.245 0.7 7.605 0.7 7.605 1.26 8.07 1.26 8.07 1.38 7.465 1.38 7.465 2.1 7.345 2.1 7.345 1.38 6.965 1.38 6.965 1.46 6.845 1.46 6.845 1.22 6.965 1.22 6.965 1.26 7.485 1.26 7.485 0.82 7.125 0.82 7.125 0.46 11.385 0.46 11.385 0.81 11.585 0.81 ;
      POLYGON 7.365 1.14 7.125 1.14 7.125 1.1 6.725 1.1 6.725 1.77 6.385 1.77 6.385 1.81 6.145 1.81 6.145 1.69 6.265 1.69 6.265 1.65 6.605 1.65 6.605 1.1 6.065 1.1 6.065 0.62 6.185 0.62 6.185 0.98 7.365 0.98 ;
      POLYGON 6.485 1.53 6.365 1.53 6.365 1.34 5.825 1.34 5.825 0.5 5.465 0.5 5.465 0.91 4.745 0.91 4.745 0.5 4.105 0.5 4.105 1.29 4.225 1.29 4.225 1.41 3.985 1.41 3.985 0.5 3.475 0.5 3.475 0.8 3.625 0.8 3.625 1.77 3.955 1.77 3.955 1.89 3.505 1.89 3.505 0.92 3.355 0.92 3.355 0.38 4.425 0.38 4.425 0.36 4.665 0.36 4.665 0.38 4.865 0.38 4.865 0.79 5.345 0.79 5.345 0.38 5.945 0.38 5.945 1.22 6.485 1.22 ;
      POLYGON 5.765 1.87 5.645 1.87 5.645 1.75 5.585 1.75 5.585 1.49 5.025 1.49 5.025 1.37 5.585 1.37 5.585 0.62 5.705 0.62 5.705 1.63 5.765 1.63 ;
      POLYGON 5.465 1.15 4.625 1.15 4.625 1.63 4.705 1.63 4.705 1.87 4.585 1.87 4.585 1.75 4.505 1.75 4.505 0.8 4.285 0.8 4.285 0.68 4.625 0.68 4.625 1.03 5.465 1.03 ;
      POLYGON 4.285 2.11 4.27 2.11 4.27 2.13 3.21 2.13 3.21 2.25 2.49 2.25 2.49 1.93 1.47 1.93 1.47 2.07 1.35 2.07 1.35 1.95 1.33 1.95 1.33 0.84 1.19 0.84 1.19 0.72 1.45 0.72 1.45 1.81 2.61 1.81 2.61 2.13 3.09 2.13 3.09 2.01 4.15 2.01 4.15 1.99 4.165 1.99 4.165 1.65 3.745 1.65 3.745 0.62 3.865 0.62 3.865 1.53 4.285 1.53 ;
      POLYGON 3.385 1.21 2.85 1.21 2.85 1.89 2.97 1.89 2.97 2.01 2.73 2.01 2.73 1.16 2.43 1.16 2.43 0.66 2.55 0.66 2.55 1.04 2.85 1.04 2.85 1.09 3.385 1.09 ;
      POLYGON 1.81 1.69 1.57 1.69 1.57 0.6 1.005 0.6 1.005 0.66 0.255 0.66 0.255 0.9 0.24 0.9 0.24 1.555 0.41 1.555 0.41 2.07 0.29 2.07 0.29 1.675 0.12 1.675 0.12 0.78 0.135 0.78 0.135 0.54 0.885 0.54 0.885 0.48 1.03 0.48 1.03 0.38 1.27 0.38 1.27 0.48 1.69 0.48 1.69 1.57 1.81 1.57 ;
  END
END SDFFX4

MACRO INVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX12 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.296 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.15 3.835 1.27 ;
        RECT 0.885 1.15 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.5 4.075 1.62 ;
        RECT 3.955 0.91 4.075 1.62 ;
        RECT 3.915 1.43 4.035 2.21 ;
        RECT 0.555 0.91 4.075 1.03 ;
        RECT 3.915 0.4 4.035 1.03 ;
        RECT 3.84 1.465 4.035 1.725 ;
        RECT 3.075 1.43 3.195 2.21 ;
        RECT 3.075 0.4 3.195 1.03 ;
        RECT 2.235 1.43 2.355 2.21 ;
        RECT 2.235 0.4 2.355 1.03 ;
        RECT 1.395 1.43 1.515 2.21 ;
        RECT 1.395 0.4 1.515 1.03 ;
        RECT 0.555 1.43 0.675 2.21 ;
        RECT 0.555 0.4 0.675 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 4.335 -0.18 4.455 0.915 ;
        RECT 3.495 -0.18 3.615 0.79 ;
        RECT 2.655 -0.18 2.775 0.79 ;
        RECT 1.815 -0.18 1.935 0.79 ;
        RECT 0.975 -0.18 1.095 0.79 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 4.335 1.43 4.455 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.43 0.255 2.79 ;
    END
  END VDD
END INVX12

MACRO DFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX8 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.645 0.725 2.965 0.845 ;
        RECT 2.665 1.34 2.785 2.085 ;
        RECT 2.645 0.725 2.765 1.46 ;
        RECT 0.265 1.025 2.765 1.145 ;
        RECT 1.945 0.665 2.065 1.46 ;
        RECT 1.825 1.34 1.945 2.085 ;
        RECT 1.105 0.665 1.225 1.46 ;
        RECT 0.985 1.34 1.105 2.08 ;
        RECT 0.265 0.885 0.51 1.145 ;
        RECT 0.265 0.665 0.385 1.46 ;
        RECT 0.145 1.34 0.265 2.08 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.885 0.86 11.125 1.04 ;
        RECT 10.745 0.885 11.005 1.09 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.414 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.41 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.0098 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.585 0.36 4.705 1.16 ;
        RECT 3.445 0.36 4.705 0.48 ;
        RECT 3.445 0.36 3.565 1.18 ;
        RECT 3.26 0.885 3.565 1.145 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.615 1.11 11.875 1.38 ;
        RECT 11.575 1.11 11.875 1.36 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.375 -0.18 11.495 0.75 ;
        RECT 10.925 0.5 11.165 0.62 ;
        RECT 10.925 -0.18 11.045 0.62 ;
        RECT 8.775 0.43 9.015 0.55 ;
        RECT 8.895 -0.18 9.015 0.55 ;
        RECT 6.395 -0.18 6.635 0.32 ;
        RECT 4.825 -0.18 4.945 0.65 ;
        RECT 3.205 -0.18 3.325 0.65 ;
        RECT 2.365 -0.18 2.485 0.655 ;
        RECT 1.525 -0.18 1.645 0.655 ;
        RECT 0.685 -0.18 0.805 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.185 1.74 11.305 2.79 ;
        RECT 9.675 2.29 9.915 2.79 ;
        RECT 8.775 2.01 8.895 2.79 ;
        RECT 8.655 2.01 8.895 2.13 ;
        RECT 6.635 2.22 6.875 2.79 ;
        RECT 5.785 2.22 6.025 2.79 ;
        RECT 4.825 1.9 5.065 2.02 ;
        RECT 4.825 1.9 4.945 2.79 ;
        RECT 3.865 1.9 4.105 2.02 ;
        RECT 3.865 1.9 3.985 2.79 ;
        RECT 3.085 1.54 3.205 2.79 ;
        RECT 2.245 1.34 2.365 2.79 ;
        RECT 1.405 1.34 1.525 2.79 ;
        RECT 0.565 1.34 0.685 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.915 0.99 11.455 0.99 11.455 1.5 11.545 1.5 11.545 1.64 11.725 1.64 11.725 1.88 11.605 1.88 11.605 1.76 11.425 1.76 11.425 1.62 11.335 1.62 11.335 1.36 10.265 1.36 10.265 1.31 10.125 1.31 10.125 1.19 10.385 1.19 10.385 1.24 11.335 1.24 11.335 0.87 11.795 0.87 11.795 0.51 11.915 0.51 ;
      POLYGON 10.665 1.99 10.545 1.99 10.545 1.6 9.885 1.6 9.885 1.56 8.695 1.56 8.695 1.15 8.815 1.15 8.815 1.44 9.885 1.44 9.885 0.6 10.125 0.6 10.125 0.72 10.005 0.72 10.005 1.48 10.665 1.48 ;
      POLYGON 10.625 1.12 10.505 1.12 10.505 0.48 9.765 0.48 9.765 1.1 9.645 1.1 9.645 0.74 9.5 0.74 9.5 0.79 8.535 0.79 8.535 0.48 7.955 0.48 7.955 0.92 7.975 0.92 7.975 1.04 7.735 1.04 7.735 0.92 7.835 0.92 7.835 0.48 7.355 0.48 7.355 1.54 6.375 1.54 6.375 1.62 6.035 1.62 6.035 0.8 5.915 0.8 5.915 0.68 6.155 0.68 6.155 1.42 7.235 1.42 7.235 0.36 8.655 0.36 8.655 0.67 9.38 0.67 9.38 0.62 9.645 0.62 9.645 0.36 10.625 0.36 ;
      POLYGON 10.445 2.25 10.205 2.25 10.205 2.17 9.015 2.17 9.015 1.89 7.935 1.89 7.935 1.21 8.335 1.21 8.335 1.33 8.055 1.33 8.055 1.77 9.135 1.77 9.135 2.05 10.325 2.05 10.325 2.13 10.445 2.13 ;
      POLYGON 10.305 1.93 9.255 1.93 9.255 1.69 9.375 1.69 9.375 1.81 10.065 1.81 10.065 1.72 10.305 1.72 ;
      POLYGON 9.405 1.32 9.285 1.32 9.285 1.03 8.575 1.03 8.575 1.65 8.175 1.65 8.175 1.53 8.455 1.53 8.455 1.03 8.175 1.03 8.175 0.6 8.415 0.6 8.415 0.91 9.405 0.91 ;
      POLYGON 8.335 2.25 7.83 2.25 7.83 2.23 7.235 2.23 7.235 2.1 5.425 2.1 5.425 2.25 5.185 2.25 5.185 2.13 5.305 2.13 5.305 1.98 7.355 1.98 7.355 2.11 7.95 2.11 7.95 2.13 8.335 2.13 ;
      POLYGON 7.715 0.72 7.595 0.72 7.595 1.99 7.475 1.99 7.475 1.86 5.665 1.86 5.665 1.78 4.065 1.78 4.065 1.04 4.185 1.04 4.185 1.66 5.665 1.66 5.665 1.26 5.645 1.26 5.645 1.02 5.785 1.02 5.785 1.74 7.475 1.74 7.475 0.6 7.715 0.6 ;
      POLYGON 7.115 1.3 6.275 1.3 6.275 1.18 6.995 1.18 6.995 0.88 7.115 0.88 ;
      POLYGON 6.855 1.06 6.615 1.06 6.615 0.56 5.705 0.56 5.705 0.9 5.425 0.9 5.425 1.4 5.545 1.4 5.545 1.54 5.305 1.54 5.305 1.4 4.585 1.4 4.585 1.54 4.345 1.54 4.345 0.92 3.945 0.92 3.945 1.42 3.625 1.42 3.625 2.08 3.505 2.08 3.505 1.42 3.02 1.42 3.02 1.2 2.885 1.2 2.885 1.08 3.14 1.08 3.14 1.3 3.825 1.3 3.825 0.72 3.925 0.72 3.925 0.6 4.045 0.6 4.045 0.8 4.465 0.8 4.465 1.28 5.305 1.28 5.305 0.78 5.585 0.78 5.585 0.44 6.735 0.44 6.735 0.94 6.855 0.94 ;
  END
END DFFRHQX8

MACRO NOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 0.99 3.335 1.11 ;
        RECT 1.695 0.99 1.935 1.13 ;
        RECT 0.65 0.99 0.8 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 1.26 2.595 1.38 ;
        RECT 2.335 1.23 2.595 1.38 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9664 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 1.5 3.575 1.62 ;
        RECT 3.455 0.73 3.575 1.62 ;
        RECT 3.205 1.23 3.575 1.38 ;
        RECT 0.555 0.73 3.575 0.85 ;
        RECT 3.075 0.61 3.195 0.85 ;
        RECT 2.555 1.5 2.675 2.21 ;
        RECT 2.235 0.61 2.355 0.85 ;
        RECT 1.395 0.61 1.515 0.85 ;
        RECT 1.275 1.5 1.395 2.21 ;
        RECT 0.555 0.61 0.675 0.85 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.435 0.48 3.675 0.6 ;
        RECT 3.435 -0.18 3.555 0.6 ;
        RECT 2.595 0.48 2.835 0.6 ;
        RECT 2.595 -0.18 2.715 0.6 ;
        RECT 1.755 0.48 1.995 0.6 ;
        RECT 1.755 -0.18 1.875 0.6 ;
        RECT 0.915 0.48 1.155 0.6 ;
        RECT 0.915 -0.18 1.035 0.6 ;
        RECT 0.135 -0.18 0.255 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.295 1.74 3.415 2.79 ;
        RECT 1.915 1.74 2.035 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
END NOR2X4

MACRO OR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X8 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.61 0.82 2.73 1.17 ;
        RECT 0.39 0.82 2.73 0.94 ;
        RECT 0.39 0.82 0.51 1.15 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.39 1.3 ;
        RECT 2.1 1.06 2.25 1.435 ;
        RECT 1.03 1.06 2.39 1.18 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.3 1.79 1.42 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.55 1.3 1.67 1.725 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 0.715 6.19 0.835 ;
        RECT 3.55 0.765 6.07 0.885 ;
        RECT 5.81 1.47 5.93 2.21 ;
        RECT 5.63 1.47 5.93 1.59 ;
        RECT 5.63 1.275 5.75 1.59 ;
        RECT 3.29 1.275 5.75 1.395 ;
        RECT 5.19 0.765 5.44 1.145 ;
        RECT 5.19 0.765 5.31 1.395 ;
        RECT 5.17 0.645 5.29 0.885 ;
        RECT 4.97 1.275 5.27 1.59 ;
        RECT 4.97 1.275 5.09 2.21 ;
        RECT 4.27 0.715 4.51 0.885 ;
        RECT 4.13 1.275 4.25 2.21 ;
        RECT 3.43 0.715 3.67 0.835 ;
        RECT 3.29 1.275 3.41 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.59 -0.18 5.71 0.645 ;
        RECT 4.75 -0.18 4.87 0.645 ;
        RECT 3.91 -0.18 4.03 0.645 ;
        RECT 2.95 0.34 3.19 0.46 ;
        RECT 2.95 -0.18 3.07 0.46 ;
        RECT 1.99 0.34 2.23 0.46 ;
        RECT 1.99 -0.18 2.11 0.46 ;
        RECT 1.03 0.34 1.27 0.46 ;
        RECT 1.03 -0.18 1.15 0.46 ;
        RECT 0.19 -0.18 0.31 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.39 1.515 5.51 2.79 ;
        RECT 4.55 1.515 4.67 2.79 ;
        RECT 3.71 1.515 3.83 2.79 ;
        RECT 2.87 1.795 2.99 2.79 ;
        RECT 0.61 1.56 0.73 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.07 1.155 2.97 1.155 2.97 1.675 1.91 1.675 1.91 2.21 1.79 2.21 1.79 1.555 2.85 1.555 2.85 0.7 0.55 0.7 0.55 0.58 2.97 0.58 2.97 1.035 5.07 1.035 ;
  END
END OR3X8

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.225 1.275 1.38 ;
        RECT 1.155 1.13 1.275 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.225 0.675 2.12 ;
        RECT 0.555 0.605 0.675 0.845 ;
        RECT 0.515 0.725 0.635 1.345 ;
        RECT 0.36 0.885 0.635 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.77 ;
        RECT 0.135 -0.18 0.255 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.5 1.095 2.79 ;
        RECT 0.135 1.47 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.74 1.395 1.74 1.395 1.01 1.035 1.01 1.035 1.105 0.755 1.105 0.755 0.985 0.915 0.985 0.915 0.89 1.395 0.89 1.395 0.53 1.515 0.53 ;
  END
END BUFX2

MACRO NOR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X8 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.605 1.205 10.985 1.325 ;
        RECT 9.585 1.23 9.845 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 1.175 8.63 1.435 ;
        RECT 8.48 1.07 8.6 1.435 ;
        RECT 6.655 1.19 8.63 1.31 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.715 1.205 5.075 1.325 ;
        RECT 3.785 1.205 4.045 1.38 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.19 2.075 1.31 ;
        RECT 1.955 1.07 2.075 1.31 ;
        RECT 1.81 1.175 1.96 1.435 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.1393 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.925 1.465 12.045 2.21 ;
        RECT 9.405 1.5 12.045 1.62 ;
        RECT 0.615 0.79 11.625 0.91 ;
        RECT 11.505 0.67 11.625 0.91 ;
        RECT 11.085 1.465 11.24 1.725 ;
        RECT 11.105 0.79 11.225 1.725 ;
        RECT 11.085 1.465 11.205 2.01 ;
        RECT 10.605 0.74 10.845 0.91 ;
        RECT 10.245 1.47 10.365 2.01 ;
        RECT 9.745 0.74 9.985 0.91 ;
        RECT 9.405 1.5 9.525 2.01 ;
        RECT 8.905 0.74 9.145 0.91 ;
        RECT 8.055 0.74 8.295 0.91 ;
        RECT 7.215 0.74 7.455 0.91 ;
        RECT 6.375 0.74 6.615 0.91 ;
        RECT 5.535 0.74 5.775 0.91 ;
        RECT 4.695 0.74 4.935 0.91 ;
        RECT 3.855 0.74 4.095 0.91 ;
        RECT 3.015 0.74 3.255 0.91 ;
        RECT 2.175 0.74 2.415 0.91 ;
        RECT 1.335 0.74 1.575 0.91 ;
        RECT 0.495 0.74 0.735 0.86 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.925 -0.18 12.045 0.67 ;
        RECT 11.085 -0.18 11.205 0.67 ;
        RECT 10.245 -0.18 10.365 0.67 ;
        RECT 9.385 -0.18 9.505 0.665 ;
        RECT 8.535 -0.18 8.655 0.67 ;
        RECT 7.695 -0.18 7.815 0.67 ;
        RECT 6.855 -0.18 6.975 0.67 ;
        RECT 6.015 -0.18 6.135 0.67 ;
        RECT 5.175 -0.18 5.295 0.67 ;
        RECT 4.335 -0.18 4.455 0.67 ;
        RECT 3.495 -0.18 3.615 0.665 ;
        RECT 2.655 -0.18 2.775 0.67 ;
        RECT 1.815 -0.18 1.935 0.67 ;
        RECT 0.975 -0.18 1.095 0.67 ;
        RECT 0.135 -0.18 0.255 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 2.655 1.795 2.775 2.79 ;
        RECT 1.815 1.795 1.935 2.79 ;
        RECT 0.975 1.795 1.095 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.625 2.25 8.985 2.25 8.985 1.675 8.265 1.675 8.265 2.01 8.145 2.01 8.145 1.675 7.395 1.675 7.395 2.01 7.275 2.01 7.275 1.675 6.555 1.675 6.555 2.01 6.435 2.01 6.435 1.465 6.555 1.465 6.555 1.555 7.275 1.555 7.275 1.465 7.395 1.465 7.395 1.555 8.145 1.555 8.145 1.47 8.265 1.47 8.265 1.555 8.985 1.555 8.985 1.47 9.105 1.47 9.105 2.13 9.825 2.13 9.825 1.74 9.945 1.74 9.945 2.13 10.665 2.13 10.665 1.74 10.785 1.74 10.785 2.13 11.505 2.13 11.505 1.74 11.625 1.74 ;
      POLYGON 8.685 2.25 6.015 2.25 6.015 1.62 5.295 1.62 5.295 2.01 5.175 2.01 5.175 1.62 4.455 1.62 4.455 2.01 4.335 2.01 4.335 1.62 3.615 1.62 3.615 2.01 3.495 2.01 3.495 1.47 3.615 1.47 3.615 1.5 4.335 1.5 4.335 1.47 4.455 1.47 4.455 1.5 5.175 1.5 5.175 1.465 5.295 1.465 5.295 1.5 6.015 1.5 6.015 1.465 6.135 1.465 6.135 2.13 6.855 2.13 6.855 1.795 6.975 1.795 6.975 2.13 7.695 2.13 7.695 1.795 7.815 1.795 7.815 2.13 8.565 2.13 8.565 1.795 8.685 1.795 ;
      POLYGON 5.715 2.25 3.075 2.25 3.075 1.675 2.355 1.675 2.355 2.21 2.235 2.21 2.235 1.675 1.515 1.675 1.515 2.21 1.395 2.21 1.395 1.675 0.675 1.675 0.675 2.21 0.555 2.21 0.555 1.465 0.675 1.465 0.675 1.555 1.395 1.555 1.395 1.465 1.515 1.465 1.515 1.555 2.235 1.555 2.235 1.47 2.355 1.47 2.355 1.555 3.075 1.555 3.075 1.47 3.195 1.47 3.195 2.13 3.915 2.13 3.915 1.74 4.035 1.74 4.035 2.13 4.755 2.13 4.755 1.74 4.875 1.74 4.875 2.13 5.595 2.13 5.595 1.74 5.715 1.74 ;
  END
END NOR4X8

MACRO AOI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.33 1.25 2.45 2.01 ;
        RECT 2.13 1.25 2.45 1.37 ;
        RECT 2.13 0.62 2.25 1.37 ;
        RECT 2.1 0.74 2.25 1.145 ;
        RECT 1.13 0.74 2.25 0.86 ;
        RECT 1.01 0.69 1.25 0.81 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.22 1.215 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.98 1.69 1.22 ;
        RECT 1.52 0.98 1.67 1.435 ;
        RECT 0.645 0.98 1.69 1.1 ;
        RECT 0.51 1.01 0.765 1.13 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.82 2.885 1.09 ;
        RECT 2.37 0.88 2.745 1.13 ;
    END
  END B0
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 1.49 1.795 1.61 2.79 ;
        RECT 0.65 1.795 0.77 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.55 -0.18 2.67 0.68 ;
        RECT 1.65 0.5 1.89 0.62 ;
        RECT 1.65 -0.18 1.77 0.62 ;
        RECT 0.43 -0.18 0.55 0.68 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.87 2.25 1.91 2.25 1.91 1.675 1.19 1.675 1.19 2.21 1.07 2.21 1.07 1.675 0.35 1.675 0.35 2.21 0.23 2.21 0.23 1.555 2.03 1.555 2.03 2.13 2.75 2.13 2.75 1.56 2.87 1.56 ;
  END
END AOI21X2

MACRO DFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX4 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.885 0.395 1.125 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.545 1.315 1.665 1.555 ;
        RECT 1.23 1.315 1.665 1.435 ;
        RECT 1.23 1.175 1.38 1.435 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.705 0.72 6.905 0.84 ;
        RECT 6.765 1.44 6.885 2.21 ;
        RECT 6.585 1.44 6.885 1.56 ;
        RECT 5.9 1.32 6.705 1.44 ;
        RECT 5.925 0.72 6.045 2.21 ;
        RECT 5.87 1.175 6.045 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.625 0.72 8.825 0.84 ;
        RECT 8.445 1.44 8.565 2.21 ;
        RECT 8.265 1.44 8.565 1.56 ;
        RECT 7.61 1.32 8.385 1.44 ;
        RECT 7.64 0.72 7.76 1.56 ;
        RECT 7.605 1.44 7.725 2.21 ;
        RECT 7.61 1.175 7.76 1.56 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.185 -0.18 9.305 0.71 ;
        RECT 8.105 -0.18 8.345 0.36 ;
        RECT 7.145 -0.18 7.385 0.36 ;
        RECT 6.185 -0.18 6.425 0.36 ;
        RECT 5.225 -0.18 5.465 0.36 ;
        RECT 4.325 -0.18 4.445 0.38 ;
        RECT 2.725 -0.18 2.845 0.38 ;
        RECT 1.485 -0.18 1.605 0.38 ;
        RECT 0.135 -0.18 0.255 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 8.865 1.58 8.985 2.79 ;
        RECT 8.025 1.56 8.145 2.79 ;
        RECT 7.185 1.56 7.305 2.79 ;
        RECT 6.345 1.56 6.465 2.79 ;
        RECT 5.505 1.56 5.625 2.79 ;
        RECT 4.605 1.67 4.725 2.79 ;
        RECT 2.825 2.26 3.065 2.79 ;
        RECT 1.385 1.95 1.505 2.79 ;
        RECT 0.135 1.46 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.725 0.9 9.545 0.9 9.545 1.46 9.405 1.46 9.405 2.21 9.285 2.21 9.285 1.46 8.725 1.46 8.725 1.22 8.845 1.22 8.845 1.34 9.425 1.34 9.425 0.78 9.605 0.78 9.605 0.66 9.725 0.66 ;
      POLYGON 9.265 1.22 9.145 1.22 9.145 0.95 8.945 0.95 8.945 0.6 5.165 0.6 5.165 1.32 5.63 1.32 5.63 1.2 5.75 1.2 5.75 1.44 5.145 1.44 5.145 2.19 5.025 2.19 5.025 1.44 4.685 1.44 4.685 1.5 4.445 1.5 4.445 1.38 4.565 1.38 4.565 1.32 5.045 1.32 5.045 0.8 4.805 0.8 4.805 0.56 4.925 0.56 4.925 0.68 5.045 0.68 5.045 0.48 9.065 0.48 9.065 0.83 9.265 0.83 ;
      POLYGON 4.925 1.16 3.945 1.16 3.945 1.89 4.085 1.89 4.085 2.01 3.825 2.01 3.825 0.84 3.685 0.84 3.685 0.72 3.945 0.72 3.945 1.04 4.925 1.04 ;
      POLYGON 4.325 2.25 3.185 2.25 3.185 2.14 2.705 2.14 2.705 2.25 1.865 2.25 1.865 1.795 1.11 1.795 1.11 1.915 1.085 1.915 1.085 2.07 0.965 2.07 0.965 1.795 0.99 1.795 0.99 0.84 0.885 0.84 0.885 0.72 1.125 0.72 1.125 0.84 1.11 0.84 1.11 1.675 1.865 1.675 1.865 1.49 1.985 1.49 1.985 2.13 2.585 2.13 2.585 2.02 3.305 2.02 3.305 2.13 4.205 2.13 4.205 1.73 4.065 1.73 4.065 1.49 4.185 1.49 4.185 1.61 4.325 1.61 ;
      POLYGON 4.085 0.5 3.965 0.5 3.965 0.54 3.565 0.54 3.565 1.42 3.705 1.42 3.705 1.66 3.585 1.66 3.585 1.54 3.445 1.54 3.445 0.54 3.085 0.54 3.085 0.62 2.465 0.62 2.465 1.66 2.345 1.66 2.345 0.6 1.845 0.6 1.845 0.62 1.245 0.62 1.245 0.6 0.675 0.6 0.675 1.58 0.555 1.58 0.555 0.48 1.045 0.48 1.045 0.38 1.365 0.38 1.365 0.5 1.725 0.5 1.725 0.48 1.805 0.48 1.805 0.38 2.045 0.38 2.045 0.48 2.465 0.48 2.465 0.5 2.965 0.5 2.965 0.42 3.845 0.42 3.845 0.38 4.085 0.38 ;
      POLYGON 3.665 2.01 3.425 2.01 3.425 1.9 3.205 1.9 3.205 1.32 2.685 1.32 2.685 1.08 2.805 1.08 2.805 1.2 3.205 1.2 3.205 0.66 3.325 0.66 3.325 1.78 3.545 1.78 3.545 1.89 3.665 1.89 ;
      POLYGON 3.085 1.69 2.965 1.69 2.965 1.9 2.345 1.9 2.345 2.01 2.105 2.01 2.105 0.84 1.965 0.84 1.965 0.72 2.225 0.72 2.225 1.78 2.845 1.78 2.845 1.57 3.085 1.57 ;
  END
END DFFX4

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.16 1.28 1.28 ;
        RECT 0.65 0.885 0.8 1.28 ;
        RECT 0.3 1.16 0.42 1.4 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 0.36 2.515 0.48 ;
        RECT 1.08 0.44 2.135 0.56 ;
        RECT 0.7 1.4 1.52 1.52 ;
        RECT 1.4 0.92 1.52 1.52 ;
        RECT 1.175 1.4 1.435 1.67 ;
        RECT 1.08 0.92 1.52 1.04 ;
        RECT 1.08 0.44 1.2 1.04 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.265 0.76 3.385 1.68 ;
        RECT 3.225 1.56 3.345 2.21 ;
        RECT 3.055 0.76 3.385 0.88 ;
        RECT 2.915 0.65 3.215 0.8 ;
        RECT 3.095 0.64 3.215 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.675 -0.18 2.795 0.69 ;
        RECT 1.655 -0.18 1.895 0.32 ;
        RECT 0.84 -0.18 0.96 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.805 1.7 2.925 2.79 ;
        RECT 0.975 2.27 1.215 2.79 ;
        RECT 0.135 1.85 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.145 1.44 3.105 1.44 3.105 1.58 2.595 1.58 2.595 2.15 0.555 2.15 0.555 1.85 0.46 1.85 0.46 1.64 0.06 1.64 0.06 0.92 0.14 0.92 0.14 0.62 0.26 0.62 0.26 1.04 0.18 1.04 0.18 1.52 0.58 1.52 0.58 1.73 0.675 1.73 0.675 2.03 2.475 2.03 2.475 1.46 2.985 1.46 2.985 1.2 3.145 1.2 ;
      POLYGON 2.865 1.34 2.355 1.34 2.355 1.62 2.145 1.62 2.145 1.74 1.905 1.74 1.905 1.62 2.025 1.62 2.025 1.5 2.235 1.5 2.235 0.8 2.135 0.8 2.135 0.68 2.375 0.68 2.375 0.8 2.355 0.8 2.355 1.22 2.865 1.22 ;
      POLYGON 2.115 1.32 1.76 1.32 1.76 1.91 1.455 1.91 1.455 1.79 1.64 1.79 1.64 0.8 1.32 0.8 1.32 0.68 1.76 0.68 1.76 1.2 2.115 1.2 ;
  END
END TBUFX1

MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 1.06 1.69 1.18 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.3 0.89 1.42 ;
        RECT 0.65 1.3 0.8 1.725 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.175 1.96 1.435 ;
        RECT 1.01 1.32 1.93 1.44 ;
        RECT 1.81 0.82 1.93 1.44 ;
        RECT 0.59 0.82 1.93 0.94 ;
        RECT 1.43 0.65 1.55 0.94 ;
        RECT 1.01 1.32 1.13 2.21 ;
        RECT 0.59 0.65 0.71 0.94 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.85 -0.18 1.97 0.7 ;
        RECT 1.01 -0.18 1.13 0.7 ;
        RECT 0.17 -0.18 0.29 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.65 1.56 1.77 2.79 ;
        RECT 0.21 1.56 0.33 2.79 ;
    END
  END VDD
END NOR2X2

MACRO TIELO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1204 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.545 0.255 0.96 ;
        RECT 0.135 0.53 0.255 0.96 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.455 1.2 0.255 1.2 0.255 1.99 0.135 1.99 0.135 1.08 0.455 1.08 ;
  END
END TIELO

MACRO SDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX1 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 1.09 0.86 1.425 ;
        RECT 0.65 1.095 0.83 1.435 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.065 0.96 6.185 1.2 ;
        RECT 5.87 0.96 6.185 1.145 ;
        RECT 5.87 0.885 6.02 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.21 7.625 1.41 ;
        RECT 7.265 1.21 7.525 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.765 0.97 7.885 1.21 ;
        RECT 7.555 0.94 7.815 1.09 ;
        RECT 6.545 0.97 7.885 1.09 ;
        RECT 6.545 0.97 6.665 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.295 0.265 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.665 -0.18 7.785 0.82 ;
        RECT 6.065 -0.18 6.185 0.64 ;
        RECT 3.795 0.39 4.035 0.51 ;
        RECT 3.795 -0.18 3.915 0.51 ;
        RECT 2.015 -0.18 2.135 0.68 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.445 1.795 7.565 2.79 ;
        RECT 6.065 1.56 6.185 2.79 ;
        RECT 3.795 2.07 4.035 2.19 ;
        RECT 3.795 2.07 3.915 2.79 ;
        RECT 1.715 2.01 1.955 2.13 ;
        RECT 1.715 2.01 1.835 2.79 ;
        RECT 0.565 1.85 0.685 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.205 0.82 8.125 0.82 8.125 1.68 8.045 1.68 8.045 1.8 7.925 1.8 7.925 1.675 6.945 1.675 6.945 1.24 7.065 1.24 7.065 1.555 8.005 1.555 8.005 0.7 8.085 0.7 8.085 0.58 8.205 0.58 ;
      POLYGON 7.145 0.85 6.425 0.85 6.425 1.56 6.825 1.56 6.825 2.21 6.705 2.21 6.705 1.68 6.305 1.68 6.305 1.44 5.355 1.44 5.355 1.59 5.255 1.59 5.255 1.99 5.135 1.99 5.135 1.47 5.235 1.47 5.235 0.72 5.135 0.72 5.135 0.6 5.375 0.6 5.375 0.72 5.355 0.72 5.355 1.32 6.305 1.32 6.305 0.73 7.025 0.73 7.025 0.59 7.145 0.59 ;
      POLYGON 5.765 1.86 5.645 1.86 5.645 1.98 5.495 1.98 5.495 2.23 4.895 2.23 4.895 0.48 4.415 0.48 4.415 0.84 4.535 0.84 4.535 1.1 4.415 1.1 4.415 0.96 4.295 0.96 4.295 0.75 3.555 0.75 3.555 0.48 3.075 0.48 3.075 0.98 3.035 0.98 3.035 1.1 3.015 1.1 3.015 1.27 2.455 1.27 2.455 1.39 2.335 1.39 2.335 1.15 2.895 1.15 2.895 0.86 2.955 0.86 2.955 0.36 3.675 0.36 3.675 0.63 4.295 0.63 4.295 0.36 5.705 0.36 5.705 0.81 5.585 0.81 5.585 0.48 5.015 0.48 5.015 1.11 5.115 1.11 5.115 1.35 5.015 1.35 5.015 2.11 5.375 2.11 5.375 1.86 5.525 1.86 5.525 1.74 5.765 1.74 ;
      POLYGON 4.775 1.99 4.655 1.99 4.655 1.56 3.755 1.56 3.755 1.13 3.875 1.13 3.875 1.44 4.655 1.44 4.655 0.72 4.535 0.72 4.535 0.6 4.775 0.6 ;
      POLYGON 4.595 2.25 4.355 2.25 4.355 1.95 3.255 1.95 3.255 2.23 2.075 2.23 2.075 1.89 1.105 1.89 1.105 2.1 0.985 2.1 0.985 1.29 1.035 1.29 1.035 0.68 1.155 0.68 1.155 1.41 1.105 1.41 1.105 1.77 2.195 1.77 2.195 2.11 3.135 2.11 3.135 1.23 3.275 1.23 3.275 1.11 3.395 1.11 3.395 1.35 3.255 1.35 3.255 1.83 4.475 1.83 4.475 2.13 4.595 2.13 ;
      POLYGON 4.195 1.32 4.055 1.32 4.055 1.01 3.635 1.01 3.635 1.59 3.495 1.59 3.495 1.71 3.375 1.71 3.375 1.47 3.515 1.47 3.515 0.99 3.195 0.99 3.195 0.6 3.435 0.6 3.435 0.87 3.635 0.87 3.635 0.89 4.175 0.89 4.175 1.08 4.195 1.08 ;
      POLYGON 2.835 0.72 2.375 0.72 2.375 1.03 2.215 1.03 2.215 1.51 2.575 1.51 2.575 1.47 2.695 1.47 2.695 1.99 2.575 1.99 2.575 1.63 1.595 1.63 1.595 1.37 1.515 1.37 1.515 1.13 1.715 1.13 1.715 1.51 2.095 1.51 2.095 0.91 2.255 0.91 2.255 0.6 2.835 0.6 ;
      POLYGON 1.975 1.39 1.855 1.39 1.855 1.01 1.395 1.01 1.395 1.53 1.475 1.53 1.475 1.65 1.235 1.65 1.235 1.53 1.275 1.53 1.275 0.56 0.915 0.56 0.915 0.97 0.52 0.97 0.52 1.24 0.4 1.24 0.4 0.85 0.795 0.85 0.795 0.44 1.715 0.44 1.715 0.89 1.975 0.89 ;
  END
END SDFFHQX1

MACRO NOR3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX4 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.18 0.97 4.42 1.09 ;
        RECT 4.18 0.82 4.3 1.09 ;
        RECT 2.84 0.82 4.3 0.94 ;
        RECT 1.86 0.97 2.96 1.09 ;
        RECT 2.84 0.82 2.96 1.09 ;
        RECT 2.045 0.94 2.305 1.09 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.92 0.99 6.16 1.2 ;
        RECT 5.815 0.93 6.075 1.16 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.63 1.08 5.4 1.2 ;
        RECT 3.72 1.21 4.75 1.33 ;
        RECT 4.63 1.08 4.75 1.33 ;
        RECT 3.72 1.06 3.84 1.33 ;
        RECT 3.08 1.06 3.84 1.18 ;
        RECT 0.94 1.21 3.2 1.33 ;
        RECT 3.08 1.06 3.2 1.33 ;
        RECT 0.94 0.885 1.09 1.33 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2416 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.58 5.66 0.7 ;
        RECT 4.2 1.69 4.32 2.21 ;
        RECT 0.36 1.69 4.32 1.81 ;
        RECT 1.64 1.69 1.76 2.21 ;
        RECT 0.36 0.58 0.48 1.81 ;
        RECT 0.07 1.465 0.48 1.585 ;
        RECT 0.07 1.465 0.22 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 5.9 -0.18 6.02 0.64 ;
        RECT 4.94 0.34 5.18 0.46 ;
        RECT 4.94 -0.18 5.06 0.46 ;
        RECT 3.98 0.34 4.22 0.46 ;
        RECT 3.98 -0.18 4.1 0.46 ;
        RECT 3.02 0.34 3.26 0.46 ;
        RECT 3.02 -0.18 3.14 0.46 ;
        RECT 2.06 0.34 2.3 0.46 ;
        RECT 2.06 -0.18 2.18 0.46 ;
        RECT 1.1 0.34 1.34 0.46 ;
        RECT 1.1 -0.18 1.22 0.46 ;
        RECT 0.14 0.34 0.38 0.46 ;
        RECT 0.14 -0.18 0.26 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 5.7 1.56 5.82 2.79 ;
        RECT 3.04 1.93 3.28 2.15 ;
        RECT 3.04 1.93 3.16 2.79 ;
        RECT 0.4 1.93 0.64 2.15 ;
        RECT 0.4 1.93 0.52 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.5 0.77 6.4 0.77 6.4 1.56 6.24 1.56 6.24 2.21 6.12 2.21 6.12 1.44 5.415 1.44 5.415 1.57 0.6 1.57 0.6 1.24 0.72 1.24 0.72 1.45 3.32 1.45 3.32 1.3 3.56 1.3 3.56 1.45 5.295 1.45 5.295 1.32 5.52 1.32 5.52 1.28 5.76 1.28 5.76 1.32 6.28 1.32 6.28 0.77 6.26 0.77 6.26 0.65 6.5 0.65 ;
  END
END NOR3BX4

MACRO INVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.79 0.415 1.245 ;
        RECT 0.295 0.76 0.415 1.245 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.125 1.515 2.015 ;
        RECT 0.65 0.76 1.515 0.88 ;
        RECT 1.395 0.59 1.515 0.88 ;
        RECT 0.65 1.125 1.515 1.245 ;
        RECT 0.65 0.76 0.8 1.245 ;
        RECT 0.65 0.71 0.77 1.485 ;
        RECT 0.555 1.365 0.675 2.015 ;
        RECT 0.555 0.59 0.675 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.365 1.095 2.79 ;
        RECT 0.135 1.365 0.255 2.79 ;
    END
  END VDD
END INVX3

MACRO CLKXOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.18 2.175 1.345 ;
        RECT 1.755 1.18 2.015 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 1.175 3.99 1.435 ;
        RECT 3.84 1.04 3.96 1.435 ;
        RECT 3.115 1.04 3.96 1.16 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 1.74 1.575 2.21 ;
        RECT 1.215 0.7 1.515 0.82 ;
        RECT 1.395 0.58 1.515 0.82 ;
        RECT 1.275 1.74 1.575 1.86 ;
        RECT 1.275 1.32 1.395 1.86 ;
        RECT 0.65 0.84 1.335 0.96 ;
        RECT 1.215 0.7 1.335 0.96 ;
        RECT 0.65 1.32 1.395 1.44 ;
        RECT 0.65 1.175 0.8 1.44 ;
        RECT 0.65 0.79 0.77 1.56 ;
        RECT 0.615 1.44 0.735 2.21 ;
        RECT 0.555 0.67 0.675 0.91 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.675 -0.18 3.795 0.68 ;
        RECT 1.815 -0.18 1.935 0.72 ;
        RECT 0.975 -0.18 1.095 0.72 ;
        RECT 0.135 -0.18 0.255 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.675 1.84 3.795 2.79 ;
        RECT 1.875 2.08 2.115 2.2 ;
        RECT 1.875 2.08 1.995 2.79 ;
        RECT 1.035 1.56 1.155 2.79 ;
        RECT 0.195 1.56 0.315 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.23 1.96 4.215 1.96 4.215 2.08 4.095 2.08 4.095 1.84 4.11 1.84 4.11 0.92 2.995 0.92 2.995 1.36 3.355 1.36 3.355 1.48 2.875 1.48 2.875 1.1 2.535 1.1 2.535 0.86 2.655 0.86 2.655 0.98 2.875 0.98 2.875 0.8 4.095 0.8 4.095 0.44 4.215 0.44 4.215 0.56 4.23 0.56 ;
      POLYGON 3.635 1.72 2.735 1.72 2.735 2.01 2.615 2.01 2.615 1.72 2.295 1.72 2.295 0.6 2.755 0.6 2.755 0.72 2.415 0.72 2.415 1.6 3.515 1.6 3.515 1.34 3.635 1.34 ;
      POLYGON 3.155 2.25 2.235 2.25 2.235 1.96 1.97 1.96 1.97 1.62 1.515 1.62 1.515 1.2 1.255 1.2 1.255 1.08 1.515 1.08 1.515 0.94 2.055 0.94 2.055 0.36 3.115 0.36 3.115 0.68 2.995 0.68 2.995 0.48 2.175 0.48 2.175 1.06 1.635 1.06 1.635 1.5 2.09 1.5 2.09 1.84 2.355 1.84 2.355 2.13 3.035 2.13 3.035 1.84 3.155 1.84 ;
  END
END CLKXOR2X4

MACRO DFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1 0 0 ;
  SIZE 10.73 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.915 1.1 2.155 1.225 ;
        RECT 1.755 1.225 2.035 1.38 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.585 1.24 7.645 1.36 ;
        RECT 6.045 1.12 6.705 1.24 ;
        RECT 6.045 0.4 6.165 1.24 ;
        RECT 5.085 0.4 6.165 0.52 ;
        RECT 3.315 1.24 5.205 1.36 ;
        RECT 5.085 0.4 5.205 1.36 ;
        RECT 4.945 0.94 5.205 1.09 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.35 1.175 9.5 1.435 ;
        RECT 9.185 1.12 9.47 1.24 ;
        RECT 9.185 1 9.305 1.24 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.335 1.015 10.66 1.15 ;
        RECT 10.51 0.885 10.66 1.15 ;
        RECT 10.335 1.015 10.455 1.26 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2744 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.5 1.495 0.74 ;
        RECT 1.365 1.585 1.485 2.03 ;
        RECT 1.23 1.465 1.435 1.725 ;
        RECT 1.315 0.62 1.435 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.73 0.18 ;
        RECT 10.475 -0.18 10.595 0.4 ;
        RECT 9.185 -0.18 9.305 0.88 ;
        RECT 7.745 -0.18 7.985 0.32 ;
        RECT 3.055 0.66 3.295 0.78 ;
        RECT 3.175 -0.18 3.295 0.78 ;
        RECT 1.795 -0.18 1.915 0.74 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.73 2.79 ;
        RECT 10.475 1.97 10.595 2.79 ;
        RECT 9.425 2.1 9.545 2.79 ;
        RECT 7.745 2.29 7.985 2.79 ;
        RECT 6.425 2.2 6.665 2.79 ;
        RECT 4.375 2.05 4.495 2.79 ;
        RECT 2.995 1.96 3.115 2.79 ;
        RECT 1.785 1.5 1.905 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.215 1.97 10.175 1.97 10.175 2.09 10.055 2.09 10.055 1.98 9.305 1.98 9.305 2.18 8.105 2.18 8.105 2.17 6.785 2.17 6.785 2.08 5.545 2.08 5.545 1.96 6.905 1.96 6.905 2.05 8.225 2.05 8.225 2.06 9.185 2.06 9.185 1.86 9.655 1.86 9.655 1.84 9.895 1.84 9.895 1.86 10.055 1.86 10.055 1.85 10.095 1.85 10.095 0.92 10.055 0.92 10.055 0.68 10.175 0.68 10.175 0.8 10.215 0.8 ;
      POLYGON 9.975 1.7 9.855 1.7 9.855 1.675 9.065 1.675 9.065 1.94 8.345 1.94 8.345 1.93 7.025 1.93 7.025 1.84 5.425 1.84 5.425 2.16 4.865 2.16 4.865 2.04 5.305 2.04 5.305 1.72 5.565 1.72 5.565 0.96 5.685 0.96 5.685 1.72 7.145 1.72 7.145 1.81 8.245 1.81 8.245 0.98 8.365 0.98 8.365 1.81 8.465 1.81 8.465 1.82 8.945 1.82 8.945 1.44 8.825 1.44 8.825 1.2 9.065 1.2 9.065 1.555 9.665 1.555 9.665 0.66 9.785 0.66 9.785 1.46 9.975 1.46 ;
      POLYGON 8.825 1.7 8.585 1.7 8.585 0.9 8.485 0.9 8.485 0.66 7.625 0.66 7.625 0.56 7.305 0.56 7.305 0.52 7.185 0.52 7.185 0.4 7.425 0.4 7.425 0.44 7.745 0.44 7.745 0.54 8.605 0.54 8.605 0.78 8.705 0.78 8.705 1.58 8.825 1.58 ;
      POLYGON 8.025 1.24 7.885 1.24 7.885 1.6 7.505 1.6 7.505 1.69 7.265 1.69 7.265 1.6 5.805 1.6 5.805 0.64 5.925 0.64 5.925 1.48 7.765 1.48 7.765 1.12 6.825 1.12 6.825 1 6.705 1 6.705 0.66 6.825 0.66 6.825 0.88 6.945 0.88 6.945 1 8.025 1 ;
      POLYGON 7.505 0.84 7.065 0.84 7.065 0.76 6.945 0.76 6.945 0.54 6.405 0.54 6.405 0.9 6.285 0.9 6.285 0.42 7.065 0.42 7.065 0.64 7.185 0.64 7.185 0.72 7.505 0.72 ;
      POLYGON 5.445 1.6 5.185 1.6 5.185 1.78 5.065 1.78 5.065 1.6 2.975 1.6 2.975 1.36 3.095 1.36 3.095 1.48 5.325 1.48 5.325 0.64 5.445 0.64 ;
      POLYGON 4.965 0.82 4.825 0.82 4.825 1.08 3.995 1.08 3.995 0.84 3.955 0.84 3.955 0.6 4.075 0.6 4.075 0.72 4.115 0.72 4.115 0.96 4.705 0.96 4.705 0.7 4.965 0.7 ;
      POLYGON 4.825 1.84 4.705 1.84 4.705 1.93 3.475 1.93 3.475 1.81 4.585 1.81 4.585 1.72 4.825 1.72 ;
      POLYGON 4.495 0.84 4.375 0.84 4.375 0.72 4.235 0.72 4.235 0.48 3.825 0.48 3.825 0.6 3.655 0.6 3.655 0.84 3.535 0.84 3.535 0.48 3.705 0.48 3.705 0.36 4.355 0.36 4.355 0.6 4.495 0.6 ;
      POLYGON 4.215 2.25 3.975 2.25 3.975 2.17 3.235 2.17 3.235 1.84 2.875 1.84 2.875 2.25 2.205 2.25 2.205 1.38 2.275 1.38 2.275 0.6 2.395 0.6 2.395 1.5 2.325 1.5 2.325 2.13 2.755 2.13 2.755 1.72 3.355 1.72 3.355 2.05 4.095 2.05 4.095 2.13 4.215 2.13 ;
      POLYGON 3.875 1.12 2.815 1.12 2.815 1.6 2.635 1.6 2.635 2.01 2.515 2.01 2.515 1.48 2.695 1.48 2.695 0.48 2.155 0.48 2.155 0.98 1.795 0.98 1.795 1.105 1.555 1.105 1.555 0.86 2.035 0.86 2.035 0.36 2.815 0.36 2.815 1 3.875 1 ;
      POLYGON 1.11 1.58 0.99 1.58 0.99 1.46 0.985 1.46 0.985 1.18 0.375 1.18 0.375 1.06 0.985 1.06 0.985 0.68 1.105 0.68 1.105 1.34 1.11 1.34 ;
  END
END DFFSRX1

MACRO AO21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.07 1.155 1.435 ;
        RECT 1.035 1.065 1.155 1.435 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.025 0.82 1.46 ;
        RECT 0.7 1 0.82 1.46 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.76 0.51 1.225 ;
        RECT 0.38 0.76 0.5 1.25 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.885 3.41 1.145 ;
        RECT 2.98 0.885 3.41 1.005 ;
        RECT 2.98 0.76 3.1 1.68 ;
        RECT 2.965 1.56 3.085 2.21 ;
        RECT 2.125 1.32 3.1 1.44 ;
        RECT 1.88 0.76 3.1 0.88 ;
        RECT 2.54 0.59 2.66 0.88 ;
        RECT 2.125 1.32 2.245 2.21 ;
        RECT 1.7 0.71 2 0.83 ;
        RECT 1.7 0.59 1.82 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 2.96 -0.18 3.08 0.64 ;
        RECT 2.12 -0.18 2.24 0.64 ;
        RECT 1.28 -0.18 1.4 0.64 ;
        RECT 0.22 -0.18 0.34 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.385 1.56 3.505 2.79 ;
        RECT 2.545 1.56 2.665 2.79 ;
        RECT 1.705 1.97 1.825 2.79 ;
        RECT 0.495 1.82 0.735 2.145 ;
        RECT 0.495 1.82 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.86 1.19 1.515 1.19 1.515 1.82 1.395 1.82 1.395 0.88 0.86 0.88 0.86 0.59 0.98 0.59 0.98 0.76 1.515 0.76 1.515 1.07 2.86 1.07 ;
      POLYGON 1.095 2.205 0.975 2.205 0.975 1.7 0.255 1.7 0.255 2.205 0.135 2.205 0.135 1.555 0.255 1.555 0.255 1.58 0.975 1.58 0.975 1.555 1.095 1.555 ;
  END
END AO21X4

MACRO SDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX2 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.71 0.885 2.83 1.44 ;
        RECT 2.68 0.885 2.83 1.26 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.74 1.16 7.885 1.4 ;
        RECT 7.61 1.175 7.785 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.585 1.17 9.965 1.36 ;
        RECT 9.585 1.165 9.845 1.38 ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.145 1.23 10.425 1.405 ;
        RECT 10.255 1.055 10.39 1.405 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.625 0.855 10.745 1.26 ;
        RECT 10.51 0.58 10.66 0.975 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.885 1.38 1.145 ;
        RECT 1.23 0.74 1.35 2.21 ;
        RECT 1.07 0.74 1.35 0.86 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.03 0.74 2.27 0.86 ;
        RECT 2.07 1.175 2.25 1.435 ;
        RECT 2.07 0.74 2.19 2.21 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.125 -0.18 10.245 0.92 ;
        RECT 7.865 -0.18 7.985 0.84 ;
        RECT 5.755 -0.18 5.995 0.38 ;
        RECT 3.875 0.64 4.115 0.76 ;
        RECT 3.995 -0.18 4.115 0.76 ;
        RECT 2.51 -0.18 2.75 0.38 ;
        RECT 1.55 -0.18 1.79 0.38 ;
        RECT 0.65 -0.18 0.77 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.965 1.62 11.085 2.79 ;
        RECT 10.065 2.1 10.185 2.79 ;
        RECT 7.765 1.84 7.885 2.79 ;
        RECT 5.715 2.2 5.835 2.79 ;
        RECT 3.875 1.98 4.115 2.1 ;
        RECT 3.875 1.98 3.995 2.79 ;
        RECT 2.49 1.56 2.61 2.79 ;
        RECT 1.65 1.58 1.77 2.79 ;
        RECT 0.81 1.56 0.93 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.985 1.5 10.665 1.5 10.665 1.98 8.825 1.98 8.825 1.72 9.105 1.72 9.105 0.84 8.985 0.84 8.985 0.6 9.105 0.6 9.105 0.72 9.225 0.72 9.225 1.86 10.545 1.86 10.545 1.38 10.865 1.38 10.865 0.68 10.985 0.68 ;
      POLYGON 9.825 0.92 9.465 0.92 9.465 1.5 9.705 1.5 9.705 1.74 9.585 1.74 9.585 1.62 9.345 1.62 9.345 0.8 9.705 0.8 9.705 0.68 9.345 0.68 9.345 0.48 8.865 0.48 8.865 0.98 8.985 0.98 8.985 1.1 8.865 1.1 8.865 1.32 8.365 1.32 8.365 1.48 8.245 1.48 8.245 1.2 8.745 1.2 8.745 0.36 9.465 0.36 9.465 0.56 9.825 0.56 ;
      POLYGON 8.625 1.08 8.125 1.08 8.125 1.6 8.525 1.6 8.525 1.96 8.405 1.96 8.405 1.72 7.175 1.72 7.175 1.78 6.895 1.78 6.895 1.66 7.055 1.66 7.055 0.68 7.175 0.68 7.175 1.6 8.005 1.6 8.005 0.96 8.505 0.96 8.505 0.6 8.625 0.6 ;
      POLYGON 7.565 0.84 7.445 0.84 7.445 0.6 7.345 0.6 7.345 0.56 6.935 0.56 6.935 1.1 6.775 1.1 6.775 1.28 6.935 1.28 6.935 1.52 6.775 1.52 6.775 1.9 7.525 1.9 7.525 2.02 6.655 2.02 6.655 0.98 6.815 0.98 6.815 0.56 6.29 0.56 6.29 0.62 5.155 0.62 5.155 1.26 5.035 1.26 5.035 0.5 6.17 0.5 6.17 0.44 6.315 0.44 6.315 0.42 6.555 0.42 6.555 0.44 7.465 0.44 7.465 0.48 7.565 0.48 ;
      POLYGON 6.695 0.86 6.535 0.86 6.535 1.84 6.415 1.84 6.415 1.44 5.535 1.44 5.535 1.32 6.415 1.32 6.415 0.74 6.695 0.74 ;
      POLYGON 6.455 2.22 6.145 2.22 6.145 2.08 5.275 2.08 5.275 2.22 5.035 2.22 5.035 2.08 4.555 2.08 4.555 1.86 2.97 1.86 2.97 0.74 3.23 0.74 3.23 0.86 3.09 0.86 3.09 1.74 4.555 1.74 4.555 1.24 4.435 1.24 4.435 1.12 4.675 1.12 4.675 1.96 6.265 1.96 6.265 2.1 6.455 2.1 ;
      POLYGON 6.115 1.2 5.415 1.2 5.415 1.72 5.355 1.72 5.355 1.84 5.235 1.84 5.235 1.6 5.295 1.6 5.295 0.86 5.275 0.86 5.275 0.74 5.515 0.74 5.515 0.86 5.415 0.86 5.415 1.08 6.115 1.08 ;
      POLYGON 4.935 1.84 4.815 1.84 4.815 1.5 4.795 1.5 4.795 0.92 4.425 0.92 4.425 1 3.895 1 3.895 1.26 3.775 1.26 3.775 0.88 4.305 0.88 4.305 0.8 4.775 0.8 4.775 0.68 4.895 0.68 4.895 0.8 4.915 0.8 4.915 1.38 4.935 1.38 ;
      POLYGON 4.315 1.44 4.135 1.44 4.135 1.5 3.635 1.5 3.635 1.62 3.395 1.62 3.395 1.5 3.515 1.5 3.515 0.62 2.51 0.62 2.51 1.24 2.37 1.24 2.37 1 2.39 1 2.39 0.62 1.91 0.62 1.91 1.46 1.79 1.46 1.79 0.62 0.39 0.62 0.39 0.52 0.27 0.52 0.27 0.4 0.51 0.4 0.51 0.5 3.635 0.5 3.635 1.38 4.015 1.38 4.015 1.32 4.315 1.32 ;
      POLYGON 1.11 1.18 0.45 1.18 0.45 1.8 0.33 1.8 0.33 0.86 0.11 0.86 0.11 0.74 0.45 0.74 0.45 1.06 1.11 1.06 ;
  END
END SDFFTRX2

MACRO SDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX2 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 1.225 1.285 1.345 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.405 1.225 0.525 1.47 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.465 1.09 1.785 ;
        RECT 0.685 1.465 1.09 1.615 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.58 ;
        RECT 2.005 1.255 2.125 1.67 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.06 0.74 7.18 1.26 ;
        RECT 7.03 0.74 7.18 1.2 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.83 1.175 8.05 1.435 ;
        RECT 7.83 0.74 7.95 2.01 ;
        RECT 7.65 0.74 7.95 0.86 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.61 0.74 8.85 0.86 ;
        RECT 8.67 0.74 8.79 2.01 ;
        RECT 8.48 0.885 8.79 1.145 ;
        RECT 8.61 0.74 8.79 1.145 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.15 -0.18 9.27 0.38 ;
        RECT 8.13 -0.18 8.37 0.38 ;
        RECT 7.17 -0.18 7.41 0.38 ;
        RECT 5.86 0.68 6.1 0.8 ;
        RECT 5.86 -0.18 5.98 0.8 ;
        RECT 4.14 -0.18 4.38 0.32 ;
        RECT 1.945 -0.18 2.065 0.86 ;
        RECT 0.545 0.68 0.785 0.8 ;
        RECT 0.545 -0.18 0.665 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.09 1.36 9.21 2.79 ;
        RECT 8.25 1.36 8.37 2.79 ;
        RECT 7.41 1.36 7.53 2.79 ;
        RECT 5.895 2.14 6.135 2.26 ;
        RECT 5.895 2.14 6.015 2.79 ;
        RECT 4.255 2.2 4.495 2.79 ;
        RECT 2.145 2.18 2.385 2.3 ;
        RECT 2.145 2.18 2.265 2.79 ;
        RECT 0.665 1.95 0.785 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.785 0.86 9.665 0.86 9.665 1.18 9.63 1.18 9.63 1.6 9.51 1.6 9.51 1.18 8.91 1.18 8.91 1.06 9.545 1.06 9.545 0.74 9.785 0.74 ;
      POLYGON 9.65 0.52 9.53 0.52 9.53 0.62 8.29 0.62 8.29 1.24 8.17 1.24 8.17 0.62 7.495 0.62 7.495 1.06 7.615 1.06 7.615 1.18 7.375 1.18 7.375 0.62 6.46 0.62 6.46 0.74 6.535 0.74 6.535 1.66 6.615 1.66 6.615 1.78 6.375 1.78 6.375 1.66 6.415 1.66 6.415 1.4 6.015 1.4 6.015 1.52 5.895 1.52 5.895 1.28 6.415 1.28 6.415 0.86 6.34 0.86 6.34 0.5 9.41 0.5 9.41 0.4 9.65 0.4 ;
      POLYGON 7.05 2.02 5.525 2.02 5.525 2.08 5.295 2.08 5.295 2.22 5.055 2.22 5.055 2.08 3.935 2.08 3.935 2.22 3.695 2.22 3.695 2.1 3.815 2.1 3.815 1.96 5.405 1.96 5.405 1.9 6.93 1.9 6.93 1.5 6.79 1.5 6.79 0.86 6.67 0.86 6.67 0.74 6.91 0.74 6.91 1.38 7.05 1.38 ;
      POLYGON 6.295 1.14 5.775 1.14 5.775 1.74 5.435 1.74 5.435 1.78 5.195 1.78 5.195 1.66 5.315 1.66 5.315 1.62 5.655 1.62 5.655 1.14 5.34 1.14 5.34 0.8 5.22 0.8 5.22 0.68 5.46 0.68 5.46 1.02 6.295 1.02 ;
      POLYGON 5.535 1.5 5.415 1.5 5.415 1.38 4.98 1.38 4.98 1.2 4.875 1.2 4.875 0.96 4.98 0.96 4.98 0.56 3.32 0.56 3.32 1.22 3.38 1.22 3.38 1.34 3.14 1.34 3.14 1.22 3.2 1.22 3.2 0.56 2.72 0.56 2.72 0.62 2.485 0.62 2.485 0.74 2.49 0.74 2.49 1.7 2.985 1.7 2.985 2.01 2.745 2.01 2.745 1.82 2.37 1.82 2.37 0.86 2.365 0.86 2.365 0.5 2.6 0.5 2.6 0.44 3.58 0.44 3.58 0.36 3.82 0.36 3.82 0.44 5.1 0.44 5.1 1.26 5.535 1.26 ;
      POLYGON 4.915 1.84 4.795 1.84 4.795 1.62 4.74 1.62 4.74 1.46 4.055 1.46 4.055 1.34 4.635 1.34 4.635 0.8 4.62 0.8 4.62 0.68 4.86 0.68 4.86 0.8 4.755 0.8 4.755 1.34 4.86 1.34 4.86 1.5 4.915 1.5 ;
      POLYGON 4.515 1.14 3.735 1.14 3.735 1.84 3.615 1.84 3.615 0.8 3.44 0.8 3.44 0.68 3.735 0.68 3.735 1.02 4.515 1.02 ;
      POLYGON 3.315 2.25 2.505 2.25 2.505 2.06 1.525 2.06 1.525 2.07 1.405 2.07 1.405 0.8 1.185 0.8 1.185 0.68 1.525 0.68 1.525 1.94 2.625 1.94 2.625 2.13 3.195 2.13 3.195 1.58 2.9 1.58 2.9 0.8 2.84 0.8 2.84 0.68 3.08 0.68 3.08 0.8 3.02 0.8 3.02 1.46 3.315 1.46 ;
      POLYGON 1.765 1.75 1.645 1.75 1.645 0.56 1.025 0.56 1.025 1.04 0.185 1.04 0.185 1.59 0.365 1.59 0.365 2.07 0.245 2.07 0.245 1.71 0.065 1.71 0.065 0.74 0.185 0.74 0.185 0.62 0.305 0.62 0.305 0.92 0.905 0.92 0.905 0.44 1.045 0.44 1.045 0.36 1.285 0.36 1.285 0.44 1.765 0.44 ;
  END
END SDFFX2

MACRO NOR3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.885 1.175 3.16 1.415 ;
        RECT 2.885 1.175 3.12 1.435 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.4 1.3 ;
        RECT 2.1 1.06 2.25 1.435 ;
        RECT 0.82 1.06 2.4 1.18 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.81 1.3 1.93 1.725 ;
        RECT 1.69 1.3 1.93 1.42 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6338 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.58 2.72 0.7 ;
        RECT 1.45 1.3 1.57 2.21 ;
        RECT 0.07 1.3 1.57 1.42 ;
        RECT 0.07 1.175 0.42 1.42 ;
        RECT 0.3 0.58 0.42 1.42 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 2.96 -0.18 3.08 0.7 ;
        RECT 2 0.34 2.24 0.46 ;
        RECT 2 -0.18 2.12 0.46 ;
        RECT 1.04 0.34 1.28 0.46 ;
        RECT 1.04 -0.18 1.16 0.46 ;
        RECT 0.08 0.34 0.32 0.46 ;
        RECT 0.08 -0.18 0.2 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 2.76 1.56 2.88 2.79 ;
        RECT 0.4 1.56 0.52 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.5 0.7 3.4 0.7 3.4 1.655 3.36 1.655 3.36 1.8 3.24 1.8 3.24 1.535 3.28 1.535 3.28 0.94 2.72 0.94 2.72 1.17 2.6 1.17 2.6 0.94 0.66 0.94 0.66 1.15 0.54 1.15 0.54 0.82 3.28 0.82 3.28 0.58 3.38 0.58 3.38 0.46 3.5 0.46 ;
  END
END NOR3BX2

MACRO AOI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X4 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.655 1.23 5.25 1.35 ;
        RECT 4.655 1.23 4.915 1.38 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.33 1.225 6.91 1.345 ;
        RECT 6.395 1.225 6.655 1.38 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.31 1.26 3.55 1.38 ;
        RECT 2.625 1.23 3.43 1.35 ;
        RECT 2.625 1.23 2.885 1.38 ;
        RECT 2.625 1.01 2.85 1.38 ;
        RECT 2.61 1.01 2.85 1.13 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 1.26 1.87 1.38 ;
        RECT 1.05 1.23 1.435 1.38 ;
        RECT 1.05 1.01 1.17 1.38 ;
        RECT 0.93 1.01 1.17 1.13 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0696 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.4 0.68 7.52 0.92 ;
        RECT 7.22 0.8 7.52 0.92 ;
        RECT 4.04 0.85 7.34 0.97 ;
        RECT 7.03 1.465 7.18 1.725 ;
        RECT 7.03 0.85 7.15 1.725 ;
        RECT 7.01 1.5 7.13 2.01 ;
        RECT 6.17 1.5 7.18 1.62 ;
        RECT 6.56 0.68 6.68 0.97 ;
        RECT 6.17 1.5 6.29 2.01 ;
        RECT 5.72 0.68 5.84 0.97 ;
        RECT 4.88 0.68 5 0.97 ;
        RECT 4.04 0.68 4.16 0.97 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 6.98 -0.18 7.1 0.73 ;
        RECT 6.14 -0.18 6.26 0.73 ;
        RECT 1.55 -0.18 1.67 0.65 ;
        RECT 0.71 -0.18 0.83 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 5.33 1.74 5.45 2.79 ;
        RECT 4.49 1.74 4.61 2.79 ;
        RECT 3.65 1.74 3.77 2.79 ;
        RECT 2.81 1.74 2.93 2.79 ;
        RECT 1.97 1.74 2.09 2.79 ;
        RECT 1.13 1.74 1.25 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.55 2.25 5.75 2.25 5.75 1.62 5.03 1.62 5.03 2.21 4.91 2.21 4.91 1.62 4.19 1.62 4.19 2.21 4.07 2.21 4.07 1.62 3.35 1.62 3.35 2.21 3.23 2.21 3.23 1.62 2.51 1.62 2.51 2.21 2.39 2.21 2.39 1.62 1.67 1.62 1.67 2.21 1.55 2.21 1.55 1.62 0.83 1.62 0.83 2.21 0.71 2.21 0.71 1.5 5.87 1.5 5.87 2.13 6.59 2.13 6.59 1.74 6.71 1.74 6.71 2.13 7.43 2.13 7.43 1.56 7.55 1.56 ;
      POLYGON 5.42 0.73 5.3 0.73 5.3 0.48 4.58 0.48 4.58 0.73 4.46 0.73 4.46 0.48 3.35 0.48 3.35 0.65 3.23 0.65 3.23 0.48 2.51 0.48 2.51 0.65 2.39 0.65 2.39 0.36 5.42 0.36 ;
      POLYGON 3.77 0.89 0.29 0.89 0.29 0.6 0.41 0.6 0.41 0.77 1.13 0.77 1.13 0.6 1.25 0.6 1.25 0.77 1.97 0.77 1.97 0.6 2.09 0.6 2.09 0.77 2.81 0.77 2.81 0.6 2.93 0.6 2.93 0.77 3.65 0.77 3.65 0.6 3.77 0.6 ;
  END
END AOI31X4

MACRO NOR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X6 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.905 1.055 7.145 1.175 ;
        RECT 6.905 0.82 7.025 1.175 ;
        RECT 4.785 0.82 7.025 0.94 ;
        RECT 3.98 1.035 4.905 1.155 ;
        RECT 4.785 0.82 4.905 1.155 ;
        RECT 4.245 1.035 4.485 1.175 ;
        RECT 3.98 0.82 4.1 1.155 ;
        RECT 2.39 0.82 4.1 0.94 ;
        RECT 2.39 0.82 2.51 1.09 ;
        RECT 1.755 0.97 2.51 1.09 ;
        RECT 1.755 0.94 2.015 1.09 ;
        RECT 1.74 1.055 1.98 1.175 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.23 7.525 1.38 ;
        RECT 6.525 1.295 7.48 1.415 ;
        RECT 7.36 1.02 7.48 1.415 ;
        RECT 5.995 1.28 6.66 1.4 ;
        RECT 5.995 1.06 6.115 1.4 ;
        RECT 5.2 1.06 6.115 1.18 ;
        RECT 5.2 1.06 5.32 1.415 ;
        RECT 4.75 1.275 5.32 1.395 ;
        RECT 3.425 1.295 4.87 1.415 ;
        RECT 3.69 1.175 3.81 1.415 ;
        RECT 3.425 1.06 3.545 1.415 ;
        RECT 2.63 1.06 3.545 1.18 ;
        RECT 2.63 1.06 2.75 1.4 ;
        RECT 2.1 1.28 2.75 1.4 ;
        RECT 1.305 1.295 2.22 1.415 ;
        RECT 1.305 1.08 1.425 1.415 ;
        RECT 0.755 1.08 1.425 1.2 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.7 1.105 7.82 1.345 ;
        RECT 7.7 1.105 7.765 1.62 ;
        RECT 0.975 1.535 7.72 1.655 ;
        RECT 7.6 1.5 7.765 1.62 ;
        RECT 7.645 1.225 7.72 1.655 ;
        RECT 5.48 1.3 5.72 1.655 ;
        RECT 2.975 1.3 3.215 1.655 ;
        RECT 0.975 1.32 1.095 1.655 ;
        RECT 0.445 1.32 1.095 1.44 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.445 1.2 0.565 1.44 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9271 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 1.775 8.06 1.895 ;
        RECT 7.94 0.58 8.06 1.895 ;
        RECT 7.9 1.465 8.06 1.895 ;
        RECT 0.555 0.58 8.06 0.7 ;
        RECT 7.28 0.4 7.4 0.9 ;
        RECT 6.96 1.775 7.08 2.21 ;
        RECT 6.32 0.4 6.44 0.7 ;
        RECT 5.36 0.4 5.48 0.7 ;
        RECT 4.585 1.775 4.705 2.21 ;
        RECT 4.4 0.4 4.52 0.915 ;
        RECT 3.44 0.4 3.56 0.7 ;
        RECT 2.48 0.4 2.6 0.7 ;
        RECT 1.84 1.775 1.96 2.21 ;
        RECT 1.515 0.4 1.635 0.915 ;
        RECT 0.555 0.4 0.675 0.92 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 6.74 0.34 6.98 0.46 ;
        RECT 6.74 -0.18 6.86 0.46 ;
        RECT 5.78 0.34 6.02 0.46 ;
        RECT 5.78 -0.18 5.9 0.46 ;
        RECT 4.82 0.34 5.06 0.46 ;
        RECT 4.82 -0.18 4.94 0.46 ;
        RECT 3.86 0.34 4.1 0.46 ;
        RECT 3.86 -0.18 3.98 0.46 ;
        RECT 2.9 0.34 3.14 0.46 ;
        RECT 2.9 -0.18 3.02 0.46 ;
        RECT 1.94 0.34 2.18 0.46 ;
        RECT 1.94 -0.18 2.06 0.46 ;
        RECT 0.975 0.34 1.215 0.46 ;
        RECT 0.975 -0.18 1.095 0.46 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.8 2.015 8.04 2.15 ;
        RECT 7.8 2.015 7.92 2.79 ;
        RECT 5.76 2.015 6 2.15 ;
        RECT 5.76 2.015 5.88 2.79 ;
        RECT 2.74 2.015 2.98 2.15 ;
        RECT 2.74 2.015 2.86 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
END NOR3X6

MACRO CLKXOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.855 1.28 0.975 1.56 ;
        RECT 0.68 1.44 0.975 1.56 ;
        RECT 0.65 1.465 0.8 1.725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 1.18 2.835 1.3 ;
        RECT 2.045 1.18 2.305 1.38 ;
        RECT 1.915 1.14 2.155 1.3 ;
        RECT 1.335 1.36 1.575 1.48 ;
        RECT 1.455 1.18 1.575 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.295 0.29 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.395 -0.18 2.515 0.78 ;
        RECT 0.495 0.55 0.735 0.67 ;
        RECT 0.615 -0.18 0.735 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.275 1.74 2.395 2.79 ;
        RECT 0.59 2.16 0.83 2.28 ;
        RECT 0.59 2.16 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.075 1.74 2.815 1.74 2.815 1.86 2.695 1.86 2.695 1.62 1.955 1.62 1.955 2.24 1.715 2.24 1.715 2.12 1.835 2.12 1.835 1.5 2.815 1.5 2.815 1.62 2.955 1.62 2.955 0.78 2.815 0.78 2.815 0.54 2.935 0.54 2.935 0.66 3.075 0.66 ;
      POLYGON 2.515 1.06 2.275 1.06 2.275 1.02 1.215 1.02 1.215 1.68 1.31 1.68 1.31 1.8 1.07 1.8 1.07 1.68 1.095 1.68 1.095 0.6 1.335 0.6 1.335 0.72 1.215 0.72 1.215 0.9 2.395 0.9 2.395 0.94 2.515 0.94 ;
      POLYGON 1.875 0.78 1.755 0.78 1.755 0.48 0.975 0.48 0.975 1.16 0.55 1.16 0.55 1.28 0.53 1.28 0.53 1.92 1.475 1.92 1.475 1.86 1.55 1.86 1.55 1.74 1.67 1.74 1.67 1.98 1.595 1.98 1.595 2.04 0.41 2.04 0.41 1.04 0.855 1.04 0.855 0.36 1.875 0.36 ;
  END
END CLKXOR2X1

MACRO NOR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X6 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.11 1.17 7.78 1.29 ;
        RECT 7.265 1.17 7.525 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.87 1.175 6.02 1.435 ;
        RECT 5.87 1.11 5.99 1.435 ;
        RECT 5.11 1.175 6.02 1.295 ;
        RECT 4.99 1.15 5.23 1.27 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.89 1.15 3.51 1.27 ;
        RECT 2.915 1.15 3.175 1.38 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.175 1.38 1.435 ;
        RECT 1.23 1.11 1.35 1.435 ;
        RECT 0.93 1.175 1.38 1.295 ;
        RECT 0.81 1.17 1.05 1.29 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.474 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.57 1.43 8.69 2.21 ;
        RECT 6.89 1.5 8.69 1.62 ;
        RECT 0.555 0.87 8.435 0.99 ;
        RECT 8.315 0.4 8.435 0.99 ;
        RECT 7.9 0.87 8.05 1.145 ;
        RECT 7.73 1.43 8.02 1.62 ;
        RECT 7.9 0.87 8.02 1.62 ;
        RECT 7.73 1.43 7.85 2.01 ;
        RECT 7.475 0.4 7.595 0.99 ;
        RECT 6.89 1.43 7.01 2.01 ;
        RECT 6.635 0.4 6.755 0.99 ;
        RECT 5.735 0.4 5.855 0.99 ;
        RECT 4.85 0.4 4.97 0.99 ;
        RECT 4.01 0.4 4.13 0.99 ;
        RECT 3.17 0.4 3.29 0.99 ;
        RECT 2.33 0.4 2.45 0.99 ;
        RECT 1.43 0.4 1.55 0.99 ;
        RECT 0.555 0.4 0.675 0.99 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.735 -0.18 8.855 0.915 ;
        RECT 7.895 -0.18 8.015 0.75 ;
        RECT 7.055 -0.18 7.175 0.75 ;
        RECT 6.155 -0.18 6.275 0.75 ;
        RECT 5.315 -0.18 5.435 0.75 ;
        RECT 4.43 -0.18 4.55 0.75 ;
        RECT 3.59 -0.18 3.71 0.75 ;
        RECT 2.75 -0.18 2.87 0.75 ;
        RECT 1.85 -0.18 1.97 0.75 ;
        RECT 1.01 -0.18 1.13 0.75 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 1.85 1.795 1.97 2.79 ;
        RECT 1.01 1.795 1.13 2.79 ;
        RECT 0.17 1.43 0.29 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.27 2.25 6.47 2.25 6.47 1.675 5.75 1.675 5.75 2.01 5.63 2.01 5.63 1.675 4.91 1.675 4.91 2.01 4.79 2.01 4.79 1.43 4.91 1.43 4.91 1.555 5.63 1.555 5.63 1.43 5.75 1.43 5.75 1.555 6.47 1.555 6.47 1.43 6.59 1.43 6.59 2.13 7.31 2.13 7.31 1.74 7.43 1.74 7.43 2.13 8.15 2.13 8.15 1.74 8.27 1.74 ;
      POLYGON 6.17 2.25 4.37 2.25 4.37 1.62 3.65 1.62 3.65 2.01 3.53 2.01 3.53 1.62 2.81 1.62 2.81 2.01 2.69 2.01 2.69 1.5 3.53 1.5 3.53 1.43 3.65 1.43 3.65 1.5 4.37 1.5 4.37 1.43 4.49 1.43 4.49 2.13 5.21 2.13 5.21 1.795 5.33 1.795 5.33 2.13 6.05 2.13 6.05 1.795 6.17 1.795 ;
      POLYGON 4.07 2.25 2.27 2.25 2.27 1.675 1.55 1.675 1.55 2.21 1.43 2.21 1.43 1.675 0.71 1.675 0.71 2.21 0.59 2.21 0.59 1.43 0.71 1.43 0.71 1.555 2.27 1.555 2.27 1.43 2.39 1.43 2.39 2.13 3.11 2.13 3.11 1.74 3.23 1.74 3.23 2.13 3.95 2.13 3.95 1.74 4.07 1.74 ;
  END
END NOR4X6

MACRO AOI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X1 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 1.175 1.12 1.45 ;
        RECT 0.85 1.205 1.035 1.46 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.3 1 2.54 1.44 ;
        RECT 2.3 1 2.42 1.46 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.94 1.2 2.18 1.44 ;
        RECT 1.81 1.175 2.07 1.435 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.885 0.51 1.44 ;
        RECT 0.36 0.885 0.51 1.355 ;
    END
  END A0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.715 1 2.86 1.345 ;
        RECT 2.66 1.085 2.835 1.435 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 1 1.68 1.46 ;
        RECT 1.52 1 1.68 1.435 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6337 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.465 3.12 1.725 ;
        RECT 2.98 0.65 3.1 1.725 ;
        RECT 1.4 0.76 3.1 0.88 ;
        RECT 2.72 0.65 3.1 0.88 ;
        RECT 2.66 1.56 3.12 1.68 ;
        RECT 2.66 1.56 2.78 2.01 ;
        RECT 1.4 0.59 1.52 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.14 -0.18 2.26 0.64 ;
        RECT 0.37 -0.18 0.49 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 1.01 1.82 1.13 2.79 ;
        RECT 0.17 1.56 0.29 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.26 2.15 3.14 2.15 3.14 2.25 1.4 2.25 1.4 1.82 1.52 1.82 1.52 2.13 2.24 2.13 2.24 1.58 2.36 1.58 2.36 2.13 3.02 2.13 3.02 1.845 3.26 1.845 ;
      POLYGON 1.94 2.01 1.82 2.01 1.82 1.7 0.71 1.7 0.71 2.21 0.59 2.21 0.59 1.56 0.71 1.56 0.71 1.58 1.82 1.58 1.82 1.56 1.94 1.56 ;
  END
END AOI222X1

MACRO SDFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX4 0 0 ;
  SIZE 14.21 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.42 0.59 1.54 2.21 ;
        RECT 0.58 1.315 1.54 1.435 ;
        RECT 0.58 1.175 0.8 1.435 ;
        RECT 0.58 0.59 0.7 2.21 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.89 0.68 4.01 2.14 ;
        RECT 2.97 1.025 4.01 1.145 ;
        RECT 3.05 0.68 3.17 2.14 ;
        RECT 2.97 0.885 3.17 1.145 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.165 0.52 8.285 0.98 ;
        RECT 7.46 0.52 8.285 0.64 ;
        RECT 7.46 0.36 7.58 0.64 ;
        RECT 5.87 0.36 7.58 0.48 ;
        RECT 5.87 0.885 6.02 1.145 ;
        RECT 5.25 1.24 5.99 1.36 ;
        RECT 5.87 0.36 5.99 1.36 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.175 1.5 11.565 1.62 ;
        RECT 11.035 1.52 11.295 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.725 1.26 11.845 1.5 ;
        RECT 11.325 1.26 11.845 1.38 ;
        RECT 11.325 1.23 11.585 1.38 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.065 1.23 13.325 1.5 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.7 1.175 13.85 1.435 ;
        RECT 13.525 1.17 13.82 1.29 ;
        RECT 13.525 0.99 13.645 1.29 ;
        RECT 12.405 0.99 13.645 1.11 ;
        RECT 12.705 0.99 12.945 1.13 ;
        RECT 12.205 1.44 12.525 1.56 ;
        RECT 12.405 0.99 12.525 1.56 ;
        RECT 12.205 1.44 12.325 1.68 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.21 0.18 ;
        RECT 13.265 -0.18 13.385 0.87 ;
        RECT 11.925 -0.18 12.045 0.63 ;
        RECT 11.025 -0.18 11.265 0.33 ;
        RECT 9.035 -0.18 9.155 0.85 ;
        RECT 7.885 -0.18 8.125 0.4 ;
        RECT 5.09 0.6 5.33 0.72 ;
        RECT 5.21 -0.18 5.33 0.72 ;
        RECT 4.31 -0.18 4.43 0.78 ;
        RECT 3.47 -0.18 3.59 0.73 ;
        RECT 2.63 -0.18 2.75 0.73 ;
        RECT 1.9 -0.18 2.02 0.53 ;
        RECT 1 -0.18 1.12 0.64 ;
        RECT 0.16 -0.18 0.28 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.21 2.79 ;
        RECT 13.185 1.9 13.305 2.79 ;
        RECT 11.725 1.9 11.845 2.79 ;
        RECT 10.915 2.17 11.035 2.79 ;
        RECT 8.745 2.29 8.985 2.79 ;
        RECT 7.545 2.12 7.785 2.24 ;
        RECT 7.545 2.12 7.665 2.79 ;
        RECT 5.99 1.96 6.23 2.08 ;
        RECT 5.99 1.96 6.11 2.79 ;
        RECT 5.15 1.72 5.27 2.79 ;
        RECT 4.31 1.62 4.43 2.79 ;
        RECT 3.47 1.49 3.59 2.79 ;
        RECT 2.63 1.49 2.75 2.79 ;
        RECT 1.84 1.97 1.96 2.79 ;
        RECT 1 1.56 1.12 2.79 ;
        RECT 0.16 1.56 0.28 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.09 1.86 13.725 1.86 13.725 2.02 13.605 2.02 13.605 1.74 12.645 1.74 12.645 1.46 12.765 1.46 12.765 1.62 13.97 1.62 13.97 0.81 13.625 0.81 13.625 0.69 14.09 0.69 ;
      POLYGON 12.805 0.81 12.35 0.81 12.35 0.87 12.085 0.87 12.085 1.8 12.485 1.8 12.485 2.04 12.365 2.04 12.365 1.92 11.965 1.92 11.965 0.87 11.685 0.87 11.685 0.57 10.785 0.57 10.785 0.48 10.215 0.48 10.215 1.21 10.165 1.21 10.165 1.75 10.045 1.75 10.045 1.09 10.095 1.09 10.095 0.36 10.905 0.36 10.905 0.45 11.805 0.45 11.805 0.75 12.23 0.75 12.23 0.69 12.805 0.69 ;
      POLYGON 11.565 0.81 11.445 0.81 11.445 0.98 10.835 0.98 10.835 1.1 10.795 1.1 10.795 1.84 11.405 1.84 11.405 1.96 10.795 1.96 10.795 2.25 10.08 2.25 10.08 2.23 9.55 2.23 9.55 2.17 7.905 2.17 7.905 2 6.74 2 6.74 1.4 6.38 1.4 6.38 1.08 6.5 1.08 6.5 1.28 6.86 1.28 6.86 1.88 8.025 1.88 8.025 2.05 9.67 2.05 9.67 2.11 10.2 2.11 10.2 2.13 10.675 2.13 10.675 0.86 11.325 0.86 11.325 0.69 11.565 0.69 ;
      POLYGON 10.665 0.72 10.555 0.72 10.555 2.01 10.435 2.01 10.435 1.99 9.805 1.99 9.805 1.93 8.145 1.93 8.145 1.76 7.3 1.76 7.3 1.24 7.22 1.24 7.22 1 7.34 1 7.34 1.12 7.42 1.12 7.42 1.64 8.265 1.64 8.265 1.81 9.805 1.81 9.805 1.45 9.765 1.45 9.765 1.17 9.885 1.17 9.885 1.33 9.925 1.33 9.925 1.87 10.435 1.87 10.435 0.72 10.425 0.72 10.425 0.6 10.665 0.6 ;
      POLYGON 9.795 0.85 9.565 0.85 9.565 1.57 9.685 1.57 9.685 1.69 9.445 1.69 9.445 1.35 8.645 1.35 8.645 1.23 9.445 1.23 9.445 0.73 9.675 0.73 9.675 0.61 9.795 0.61 ;
      POLYGON 9.225 1.11 8.525 1.11 8.525 1.57 8.625 1.57 8.625 1.69 8.385 1.69 8.385 1.57 8.405 1.57 8.405 1.22 7.76 1.22 7.76 1.4 7.88 1.4 7.88 1.52 7.64 1.52 7.64 0.88 6.94 0.88 6.94 0.72 6.82 0.72 6.82 0.6 7.06 0.6 7.06 0.76 7.76 0.76 7.76 1.1 8.405 1.1 8.405 0.99 8.645 0.99 8.645 0.4 8.765 0.4 8.765 0.99 9.225 0.99 ;
      POLYGON 7.18 1.6 7.06 1.6 7.06 1.48 6.98 1.48 6.98 1.16 6.7 1.16 6.7 0.96 6.26 0.96 6.26 1.6 5.01 1.6 5.01 1.54 4.97 1.54 4.97 1.3 5.09 1.3 5.09 1.42 5.13 1.42 5.13 1.48 6.14 1.48 6.14 0.84 6.4 0.84 6.4 0.6 6.64 0.6 6.64 0.72 6.52 0.72 6.52 0.84 6.82 0.84 6.82 1.04 7.1 1.04 7.1 1.36 7.18 1.36 ;
      POLYGON 6.62 1.64 6.5 1.64 6.5 1.84 5.81 1.84 5.81 1.96 5.57 1.96 5.57 1.84 5.69 1.84 5.69 1.72 6.38 1.72 6.38 1.52 6.62 1.52 ;
      POLYGON 5.75 1.12 4.85 1.12 4.85 2.14 4.73 2.14 4.73 1.12 4.29 1.12 4.29 1.24 4.17 1.24 4.17 1 4.73 1 4.73 0.64 4.85 0.64 4.85 1 5.63 1 5.63 0.88 5.75 0.88 ;
      POLYGON 2.33 1.82 2.21 1.82 2.21 1.42 1.66 1.42 1.66 1.3 2.21 1.3 2.21 0.68 2.33 0.68 ;
  END
END SDFFSX4

MACRO DFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX8 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.79 0.655 2.91 2.21 ;
        RECT 0.07 1.025 2.91 1.145 ;
        RECT 1.95 0.655 2.07 2.21 ;
        RECT 1.11 0.655 1.23 2.205 ;
        RECT 0.27 0.655 0.39 2.205 ;
        RECT 0.07 0.885 0.39 1.145 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.84 0.49 7.96 1.23 ;
        RECT 7.34 0.49 7.96 0.61 ;
        RECT 7.34 0.36 7.46 0.61 ;
        RECT 5.58 0.36 7.46 0.48 ;
        RECT 5.58 0.885 5.73 1.145 ;
        RECT 5.58 0.36 5.7 1.34 ;
        RECT 5.16 1.22 5.7 1.34 ;
        RECT 5.04 1.26 5.28 1.38 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.16 1.14 10.425 1.385 ;
        RECT 10.165 1.12 10.425 1.385 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.6 1.21 11.005 1.385 ;
        RECT 10.745 1.18 11.005 1.385 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.4 -0.18 10.52 0.74 ;
        RECT 8.82 0.46 9.06 0.58 ;
        RECT 8.82 -0.18 8.94 0.58 ;
        RECT 7.58 -0.18 7.82 0.37 ;
        RECT 4.84 -0.18 4.96 0.68 ;
        RECT 4 -0.18 4.12 0.73 ;
        RECT 3.27 -0.18 3.39 0.53 ;
        RECT 2.37 -0.18 2.49 0.645 ;
        RECT 1.53 -0.18 1.65 0.645 ;
        RECT 0.69 -0.18 0.81 0.645 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.28 1.745 10.4 2.79 ;
        RECT 8.88 2.07 9 2.79 ;
        RECT 8.76 2.07 9 2.19 ;
        RECT 8.16 2.29 8.4 2.79 ;
        RECT 5.62 1.98 5.86 2.15 ;
        RECT 5.62 1.98 5.74 2.79 ;
        RECT 4.84 1.74 4.96 2.79 ;
        RECT 4 1.56 4.12 2.79 ;
        RECT 3.21 1.97 3.33 2.79 ;
        RECT 2.37 1.465 2.49 2.79 ;
        RECT 1.53 1.465 1.65 2.79 ;
        RECT 0.69 1.465 0.81 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.94 0.74 10.76 0.74 10.76 1 10.04 1 10.04 1.505 10.82 1.505 10.82 1.9 10.7 1.9 10.7 1.625 10.04 1.625 10.04 2.23 9.56 2.23 9.56 2.25 9.32 2.25 9.32 2.13 9.36 2.13 9.36 1.95 8.64 1.95 8.64 2.07 8.375 2.07 8.375 2.17 8.04 2.17 8.04 2.25 7.48 2.25 7.48 2.13 7.92 2.13 7.92 2.05 8.255 2.05 8.255 1.95 8.52 1.95 8.52 1.83 9.48 1.83 9.48 2.11 9.92 2.11 9.92 1 9.84 1 9.84 0.88 10.64 0.88 10.64 0.62 10.82 0.62 10.82 0.5 10.94 0.5 ;
      POLYGON 9.74 0.76 9.72 0.76 9.72 1.99 9.6 1.99 9.6 1.33 8.56 1.33 8.56 1.21 9.6 1.21 9.6 0.64 9.62 0.64 9.62 0.5 9.74 0.5 ;
      POLYGON 9.48 1.08 9.36 1.08 9.36 0.84 8.58 0.84 8.58 0.55 8.2 0.55 8.2 1.47 7.44 1.47 7.44 1.65 7.56 1.65 7.56 1.77 7.32 1.77 7.32 0.9 6.62 0.9 6.62 0.66 6.74 0.66 6.74 0.78 7.1 0.78 7.1 0.73 7.34 0.73 7.34 0.78 7.44 0.78 7.44 1.35 8.08 1.35 8.08 0.43 8.7 0.43 8.7 0.72 9.48 0.72 ;
      POLYGON 9.22 1.09 8.44 1.09 8.44 1.47 8.46 1.47 8.46 1.71 8.4 1.71 8.4 1.83 7.8 1.83 7.8 2.01 7.11 2.01 7.11 2.21 6.99 2.21 6.99 1.69 7.01 1.69 7.01 1.14 6.38 1.14 6.38 0.72 6.24 0.72 6.24 0.6 6.5 0.6 6.5 1.02 7.13 1.02 7.13 1.89 7.68 1.89 7.68 1.71 8.28 1.71 8.28 1.59 8.32 1.59 8.32 0.79 8.34 0.79 8.34 0.67 8.46 0.67 8.46 0.97 9.22 0.97 ;
      POLYGON 6.89 1.38 6.09 1.38 6.09 1.1 6.21 1.1 6.21 1.26 6.89 1.26 ;
      POLYGON 6.69 2.21 6.57 2.21 6.57 1.62 4.8 1.62 4.8 1.42 4.64 1.42 4.64 1.3 4.92 1.3 4.92 1.5 5.85 1.5 5.85 0.72 5.82 0.72 5.82 0.6 6.06 0.6 6.06 0.72 5.97 0.72 5.97 1.5 6.69 1.5 ;
      POLYGON 6.27 2.21 6.15 2.21 6.15 1.86 5.38 1.86 5.38 2.21 5.26 2.21 5.26 1.74 6.27 1.74 ;
      POLYGON 5.46 1.1 4.52 1.1 4.52 1.56 4.54 1.56 4.54 2.21 4.42 2.21 4.42 1.68 4.4 1.68 4.4 1.1 3.7 1.1 3.7 1.82 3.58 1.82 3.58 1.1 3.19 1.1 3.19 1.22 3.07 1.22 3.07 0.98 3.58 0.98 3.58 0.68 3.7 0.68 3.7 0.98 4.4 0.98 4.4 0.86 4.42 0.86 4.42 0.63 4.54 0.63 4.54 0.98 5.34 0.98 5.34 0.86 5.46 0.86 ;
  END
END DFFSHQX8

MACRO NOR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X4 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.055 0.97 4.295 1.09 ;
        RECT 4.055 0.82 4.175 1.09 ;
        RECT 1.855 0.82 4.175 0.94 ;
        RECT 1.735 0.97 2.015 1.09 ;
        RECT 1.755 0.94 2.015 1.09 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.875 1.01 4.995 1.25 ;
        RECT 4.71 1.01 4.995 1.145 ;
        RECT 4.71 0.885 4.86 1.145 ;
        RECT 3.595 1.21 4.73 1.33 ;
        RECT 4.61 1.025 4.73 1.33 ;
        RECT 3.595 1.06 3.715 1.33 ;
        RECT 2.8 1.06 3.715 1.18 ;
        RECT 2.255 1.07 2.92 1.19 ;
        RECT 1.475 1.21 2.39 1.33 ;
        RECT 2.255 1.07 2.39 1.33 ;
        RECT 1.475 1.08 1.595 1.33 ;
        RECT 0.975 1.08 1.595 1.2 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 1.45 5.335 1.57 ;
        RECT 5.215 1.24 5.335 1.57 ;
        RECT 3.095 1.3 3.335 1.57 ;
        RECT 0.92 1.32 1.04 1.57 ;
        RECT 0.39 1.32 1.04 1.44 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2416 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.455 1.465 5.73 1.725 ;
        RECT 1.835 1.69 5.575 1.81 ;
        RECT 5.455 0.58 5.575 1.81 ;
        RECT 0.495 0.58 5.575 0.7 ;
        RECT 4.395 1.69 4.515 2.21 ;
        RECT 1.835 1.69 1.955 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.775 0.34 6.015 0.46 ;
        RECT 5.775 -0.18 5.895 0.46 ;
        RECT 4.815 0.34 5.055 0.46 ;
        RECT 4.815 -0.18 4.935 0.46 ;
        RECT 3.855 0.34 4.095 0.46 ;
        RECT 3.855 -0.18 3.975 0.46 ;
        RECT 2.895 0.34 3.135 0.46 ;
        RECT 2.895 -0.18 3.015 0.46 ;
        RECT 1.935 0.34 2.175 0.46 ;
        RECT 1.935 -0.18 2.055 0.46 ;
        RECT 0.975 0.34 1.215 0.46 ;
        RECT 0.975 -0.18 1.095 0.46 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.295 1.93 5.535 2.15 ;
        RECT 5.295 1.93 5.415 2.79 ;
        RECT 2.955 1.93 3.195 2.15 ;
        RECT 2.955 1.93 3.075 2.79 ;
        RECT 0.555 1.56 0.675 2.79 ;
    END
  END VDD
END NOR3X4

MACRO CLKINVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX3 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.79 0.415 1.245 ;
        RECT 0.295 0.76 0.415 1.245 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.125 1.515 2.015 ;
        RECT 0.65 0.76 1.515 0.88 ;
        RECT 1.395 0.59 1.515 0.88 ;
        RECT 0.65 1.125 1.515 1.245 ;
        RECT 0.65 0.76 0.8 1.245 ;
        RECT 0.65 0.71 0.77 1.485 ;
        RECT 0.555 1.365 0.675 2.015 ;
        RECT 0.555 0.59 0.675 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.365 1.095 2.79 ;
        RECT 0.135 1.365 0.255 2.79 ;
    END
  END VDD
END CLKINVX3

MACRO SDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX4 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.185 0.63 2.305 0.87 ;
        RECT 1.965 1.315 2.205 1.65 ;
        RECT 2.085 0.75 2.205 1.65 ;
        RECT 1.23 1.315 2.205 1.435 ;
        RECT 1.345 0.63 1.465 0.87 ;
        RECT 1.005 1.53 1.38 1.65 ;
        RECT 1.23 1.175 1.38 1.65 ;
        RECT 1.26 0.75 1.38 1.65 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.685 1.295 ;
        RECT 0.565 1.055 0.685 1.295 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.595 1.2 7.715 1.44 ;
        RECT 7.32 1.315 7.715 1.435 ;
        RECT 7.32 1.175 7.47 1.435 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.715 1.23 9.06 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.005 0.99 9.375 1.11 ;
        RECT 8.235 0.97 9.265 1.09 ;
        RECT 9.005 0.94 9.265 1.11 ;
        RECT 8.075 1.19 8.355 1.31 ;
        RECT 8.235 0.97 8.355 1.31 ;
        RECT 8.075 1.19 8.195 1.44 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.135 -0.18 9.255 0.82 ;
        RECT 7.755 -0.18 7.875 0.83 ;
        RECT 5.465 0.39 5.705 0.51 ;
        RECT 5.585 -0.18 5.705 0.51 ;
        RECT 3.445 -0.18 3.565 0.68 ;
        RECT 2.605 -0.18 2.725 0.68 ;
        RECT 1.765 -0.18 1.885 0.68 ;
        RECT 0.925 -0.18 1.045 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 8.975 1.795 9.095 2.79 ;
        RECT 7.595 1.85 7.715 2.79 ;
        RECT 5.465 2.07 5.705 2.19 ;
        RECT 5.465 2.07 5.585 2.79 ;
        RECT 3.405 2.01 3.645 2.13 ;
        RECT 3.405 2.01 3.525 2.79 ;
        RECT 2.445 2.01 2.685 2.13 ;
        RECT 2.445 2.01 2.565 2.79 ;
        RECT 1.485 2.01 1.725 2.13 ;
        RECT 1.485 2.01 1.605 2.79 ;
        RECT 0.585 2.11 0.705 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.675 0.82 9.615 0.82 9.615 1.68 9.575 1.68 9.575 1.8 9.455 1.8 9.455 1.675 8.475 1.675 8.475 1.24 8.595 1.24 8.595 1.555 9.495 1.555 9.495 0.7 9.555 0.7 9.555 0.58 9.675 0.58 ;
      POLYGON 8.615 0.85 8.115 0.85 8.115 1.07 7.955 1.07 7.955 1.56 8.355 1.56 8.355 2.21 8.235 2.21 8.235 1.68 7.025 1.68 7.025 1.76 6.785 1.76 6.785 1.53 6.905 1.53 6.905 0.72 6.885 0.72 6.885 0.6 7.125 0.6 7.125 0.72 7.025 0.72 7.025 1.56 7.835 1.56 7.835 0.95 7.995 0.95 7.995 0.73 8.495 0.73 8.495 0.59 8.615 0.59 ;
      POLYGON 7.455 0.83 7.335 0.83 7.335 0.48 6.765 0.48 6.765 1.39 6.665 1.39 6.665 1.88 7.235 1.88 7.235 2.03 7.355 2.03 7.355 2.15 7.115 2.15 7.115 2 6.545 2 6.545 1.15 6.645 1.15 6.645 0.48 6.165 0.48 6.165 0.88 6.185 0.88 6.185 1.12 6.045 1.12 6.045 0.75 5.225 0.75 5.225 0.48 4.745 0.48 4.745 1 4.665 1 4.665 1.25 4.125 1.25 4.125 1.37 4.005 1.37 4.005 1.13 4.545 1.13 4.545 0.88 4.625 0.88 4.625 0.36 5.345 0.36 5.345 0.63 6.045 0.63 6.045 0.36 7.455 0.36 ;
      POLYGON 6.525 0.72 6.425 0.72 6.425 1.99 6.305 1.99 6.305 1.36 5.485 1.36 5.485 1.31 5.365 1.31 5.365 1.19 5.605 1.19 5.605 1.24 6.305 1.24 6.305 0.72 6.285 0.72 6.285 0.6 6.525 0.6 ;
      POLYGON 6.265 2.25 6.025 2.25 6.025 1.95 4.925 1.95 4.925 2.23 3.845 2.23 3.845 1.89 0.135 1.89 0.135 1.675 0.12 1.675 0.12 0.935 0.325 0.935 0.325 0.63 0.445 0.63 0.445 1.055 0.24 1.055 0.24 1.555 0.255 1.555 0.255 1.77 3.965 1.77 3.965 2.11 4.805 2.11 4.805 1.23 4.885 1.23 4.885 1.11 5.005 1.11 5.005 1.35 4.925 1.35 4.925 1.83 6.145 1.83 6.145 2.13 6.265 2.13 ;
      POLYGON 5.925 1.07 5.245 1.07 5.245 1.59 5.165 1.59 5.165 1.71 5.045 1.71 5.045 1.47 5.125 1.47 5.125 0.99 4.865 0.99 4.865 0.6 5.105 0.6 5.105 0.87 5.245 0.87 5.245 0.95 5.925 0.95 ;
      POLYGON 4.505 0.72 3.885 0.72 3.885 1.49 4.245 1.49 4.245 1.47 4.365 1.47 4.365 1.99 4.245 1.99 4.245 1.61 3.765 1.61 3.765 1.37 3.185 1.37 3.185 1.13 3.305 1.13 3.305 1.25 3.765 1.25 3.765 0.6 4.505 0.6 ;
      POLYGON 3.645 1.13 3.525 1.13 3.525 1.01 3.065 1.01 3.065 1.53 3.165 1.53 3.165 1.65 2.925 1.65 2.925 1.53 2.945 1.53 2.945 1.01 2.545 1.01 2.545 1.19 2.425 1.19 2.425 0.89 2.945 0.89 2.945 0.66 3.025 0.66 3.025 0.54 3.145 0.54 3.145 0.89 3.645 0.89 ;
  END
END SDFFHQX4

MACRO OAI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X2 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.035 1.06 4.535 1.18 ;
        RECT 3.26 1.06 3.41 1.435 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.555 0.82 2.675 1.15 ;
        RECT 2.39 0.82 2.675 1.145 ;
        RECT 0.595 0.82 2.675 0.94 ;
        RECT 0.595 0.82 0.715 1.15 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.53 1.3 3.77 1.42 ;
        RECT 3.55 1.3 3.7 1.725 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.27 1.3 ;
        RECT 2.1 1.06 2.25 1.435 ;
        RECT 0.975 1.06 2.27 1.18 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.3 1.57 1.42 ;
        RECT 1.23 1.465 1.38 1.725 ;
        RECT 1.26 1.3 1.38 1.725 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.215 0.65 4.455 0.77 ;
        RECT 3.375 0.76 4.335 0.88 ;
        RECT 3.575 1.845 3.695 2.21 ;
        RECT 3.375 0.65 3.615 0.88 ;
        RECT 2.795 1.845 3.695 1.965 ;
        RECT 2.795 0.82 3.495 0.94 ;
        RECT 2.795 0.82 2.915 1.965 ;
        RECT 1.67 1.56 2.915 1.68 ;
        RECT 2.625 1.52 2.915 1.68 ;
        RECT 1.67 1.56 1.79 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 2.475 0.34 2.715 0.46 ;
        RECT 2.475 -0.18 2.595 0.46 ;
        RECT 1.515 0.34 1.755 0.46 ;
        RECT 1.515 -0.18 1.635 0.46 ;
        RECT 0.555 0.34 0.795 0.46 ;
        RECT 0.555 -0.18 0.675 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.215 1.56 4.335 2.79 ;
        RECT 2.815 2.085 3.055 2.205 ;
        RECT 2.815 2.085 2.935 2.79 ;
        RECT 0.555 1.56 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.815 0.65 4.695 0.65 4.695 0.53 3.975 0.53 3.975 0.64 3.855 0.64 3.855 0.53 3.135 0.53 3.135 0.7 0.075 0.7 0.075 0.58 3.015 0.58 3.015 0.41 3.855 0.41 3.855 0.4 3.975 0.4 3.975 0.41 4.815 0.41 ;
  END
END OAI32X2

MACRO TLATNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX1 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.4 0.76 1.52 ;
        RECT 0.64 1.02 0.76 1.52 ;
        RECT 0.36 1.05 0.51 1.52 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.195 1.165 3.465 1.38 ;
        RECT 3.195 1.09 3.315 1.47 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 1.175 3.99 1.435 ;
        RECT 3.855 0.68 3.975 2.15 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.085 0.68 5.205 2.12 ;
        RECT 4.945 0.94 5.205 1.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.665 -0.18 4.785 0.73 ;
        RECT 3.435 -0.18 3.555 0.73 ;
        RECT 1.86 -0.18 1.98 0.64 ;
        RECT 0.58 -0.18 0.7 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.665 1.47 4.785 2.79 ;
        RECT 3.435 1.5 3.555 2.79 ;
        RECT 2.06 2.23 2.18 2.79 ;
        RECT 0.62 1.88 0.74 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.965 1.33 4.365 1.33 4.365 2.12 4.245 2.12 4.245 0.68 4.365 0.68 4.365 1.21 4.965 1.21 ;
      POLYGON 3.705 1.24 3.585 1.24 3.585 0.97 3.195 0.97 3.195 0.56 2.52 0.56 2.52 1.63 2.66 1.63 2.66 1.87 2.54 1.87 2.54 1.75 2.4 1.75 2.4 1.35 2.04 1.35 2.04 1.47 1.92 1.47 1.92 1.23 2.4 1.23 2.4 0.64 2.28 0.64 2.28 0.4 2.4 0.4 2.4 0.44 3.315 0.44 3.315 0.85 3.705 0.85 ;
      POLYGON 3.075 2.11 1.75 2.11 1.75 2.15 1.12 2.15 1.12 1.43 1.38 1.43 1.38 0.9 0.36 0.9 0.36 0.78 1.5 0.78 1.5 1.31 1.56 1.31 1.56 1.55 1.24 1.55 1.24 2.03 1.63 2.03 1.63 1.99 2.955 1.99 2.955 0.68 3.075 0.68 ;
      POLYGON 2.28 1.06 1.8 1.06 1.8 1.79 1.48 1.79 1.48 1.91 1.36 1.91 1.36 1.67 1.68 1.67 1.68 1.06 1.62 1.06 1.62 0.64 1.22 0.64 1.22 0.4 1.34 0.4 1.34 0.52 1.74 0.52 1.74 0.94 2.16 0.94 2.16 0.82 2.28 0.82 ;
      POLYGON 1.26 1.22 1 1.22 1 1.76 0.26 1.76 0.26 1.88 0.14 1.88 0.14 1.76 0.12 1.76 0.12 0.52 0.16 0.52 0.16 0.4 0.28 0.4 0.28 0.64 0.24 0.64 0.24 1.64 0.88 1.64 0.88 1.1 1.26 1.1 ;
  END
END TLATNX1

MACRO AO21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X2 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 1 1.38 1.46 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 0.99 0.955 1.23 ;
        RECT 0.65 0.99 0.955 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.065 0.51 1.52 ;
        RECT 0.39 0.95 0.51 1.52 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.225 1.295 2.345 2.21 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.975 1.055 2.22 1.175 ;
        RECT 1.975 0.59 2.095 1.175 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 2.395 -0.18 2.515 0.64 ;
        RECT 1.555 -0.18 1.675 0.64 ;
        RECT 0.335 -0.18 0.455 0.83 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.645 1.56 2.765 2.79 ;
        RECT 1.805 1.97 1.925 2.79 ;
        RECT 0.615 2.1 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.855 1.23 1.62 1.23 1.62 1.7 1.615 1.7 1.615 1.82 1.495 1.82 1.495 1.58 1.5 1.58 1.5 0.88 1.075 0.88 1.075 0.59 1.195 0.59 1.195 0.76 1.62 0.76 1.62 0.99 1.855 0.99 ;
      RECT 0.075 1.64 1.255 1.76 ;
  END
END AO21X2

MACRO AOI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.76 3.41 1.21 ;
        RECT 3.26 0.76 3.38 1.235 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.32 0.885 2.54 1.145 ;
        RECT 2.32 0.75 2.51 1.145 ;
        RECT 2.32 0.75 2.44 1.15 ;
        RECT 0.48 0.75 2.51 0.87 ;
        RECT 0.48 0.75 0.6 1.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 0.99 2.16 1.11 ;
        RECT 0.94 0.99 1.09 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.23 1.725 1.5 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.08 1.355 3.2 2.01 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 3 0.4 3.12 1.475 ;
        RECT 1.44 0.51 3.12 0.63 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.42 -0.18 3.54 0.64 ;
        RECT 2.46 -0.18 2.7 0.39 ;
        RECT 0.28 0.46 0.52 0.58 ;
        RECT 0.28 -0.18 0.4 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 2.24 1.86 2.36 2.79 ;
        RECT 1.4 1.86 1.52 2.79 ;
        RECT 0.56 1.86 0.68 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.62 2.25 2.66 2.25 2.66 1.74 1.94 1.74 1.94 2.21 1.82 2.21 1.82 1.74 1.1 1.74 1.1 2.21 0.98 2.21 0.98 1.74 0.26 1.74 0.26 2.21 0.14 2.21 0.14 1.56 0.26 1.56 0.26 1.62 0.98 1.62 0.98 1.56 1.1 1.56 1.1 1.62 2.66 1.62 2.66 1.56 2.78 1.56 2.78 2.13 3.5 2.13 3.5 1.56 3.62 1.56 ;
  END
END AOI31X2

MACRO NOR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.555 0.82 2.675 1.15 ;
        RECT 0.39 0.82 2.675 0.94 ;
        RECT 0.39 0.82 0.51 1.15 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.335 1.3 ;
        RECT 2.1 1.06 2.25 1.435 ;
        RECT 0.975 1.06 2.335 1.18 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.605 1.3 1.845 1.42 ;
        RECT 1.465 1.52 1.725 1.67 ;
        RECT 1.605 1.3 1.725 1.67 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6208 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.795 0.595 3.12 0.855 ;
        RECT 1.735 1.79 2.915 1.91 ;
        RECT 2.795 0.58 2.915 1.91 ;
        RECT 0.495 0.58 2.915 0.7 ;
        RECT 1.735 1.79 1.855 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.895 0.34 3.135 0.46 ;
        RECT 2.895 -0.18 3.015 0.46 ;
        RECT 1.935 0.34 2.175 0.46 ;
        RECT 1.935 -0.18 2.055 0.46 ;
        RECT 0.975 0.34 1.215 0.46 ;
        RECT 0.975 -0.18 1.095 0.46 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.635 2.03 2.875 2.15 ;
        RECT 2.635 2.03 2.755 2.79 ;
        RECT 0.555 1.56 0.675 2.79 ;
    END
  END VDD
END NOR3X2

MACRO NAND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X8 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.605 1.03 10.97 1.15 ;
        RECT 9.585 0.94 9.845 1.09 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.9 1.175 8.05 1.435 ;
        RECT 7.865 1.055 7.985 1.295 ;
        RECT 6.655 1.175 8.05 1.295 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.775 1.175 5.075 1.295 ;
        RECT 3.84 1.175 3.99 1.435 ;
        RECT 3.775 1.055 3.895 1.295 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.175 2.075 1.295 ;
        RECT 1.955 1.055 2.075 1.295 ;
        RECT 1.81 1.175 1.96 1.435 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.9616 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.345 0.7 12.105 0.82 ;
        RECT 11.505 1.47 11.625 2.21 ;
        RECT 0.555 1.555 11.625 1.675 ;
        RECT 11.09 0.7 11.24 1.145 ;
        RECT 11.09 0.7 11.21 1.675 ;
        RECT 10.645 1.47 10.765 2.21 ;
        RECT 9.805 1.465 9.925 2.21 ;
        RECT 8.965 1.47 9.085 2.21 ;
        RECT 8.115 1.555 8.235 2.21 ;
        RECT 7.275 1.465 7.395 2.21 ;
        RECT 6.435 1.465 6.555 2.21 ;
        RECT 5.595 1.47 5.715 2.21 ;
        RECT 4.755 1.47 4.875 2.21 ;
        RECT 3.915 1.555 4.035 2.21 ;
        RECT 3.075 1.47 3.195 2.21 ;
        RECT 2.235 1.555 2.355 2.21 ;
        RECT 1.395 1.465 1.515 2.21 ;
        RECT 0.555 1.465 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 2.655 -0.18 2.775 0.645 ;
        RECT 1.815 -0.18 1.935 0.645 ;
        RECT 0.975 -0.18 1.095 0.645 ;
        RECT 0.135 -0.18 0.255 0.645 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.925 1.47 12.045 2.79 ;
        RECT 11.085 1.795 11.205 2.79 ;
        RECT 10.225 1.795 10.345 2.79 ;
        RECT 9.385 1.795 9.505 2.79 ;
        RECT 8.535 1.795 8.655 2.79 ;
        RECT 7.695 1.795 7.815 2.79 ;
        RECT 6.855 1.795 6.975 2.79 ;
        RECT 6.015 1.795 6.135 2.79 ;
        RECT 5.175 1.795 5.295 2.79 ;
        RECT 4.335 1.795 4.455 2.79 ;
        RECT 3.495 1.795 3.615 2.79 ;
        RECT 2.655 1.795 2.775 2.79 ;
        RECT 1.815 1.795 1.935 2.79 ;
        RECT 0.975 1.795 1.095 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      RECT 6.375 0.46 11.685 0.58 ;
      POLYGON 8.745 0.82 6.015 0.82 6.015 0.595 3.435 0.595 3.435 0.475 6.135 0.475 6.135 0.7 8.745 0.7 ;
      POLYGON 5.775 0.835 5.655 0.835 5.655 0.885 0.615 0.885 0.615 0.84 0.495 0.84 0.495 0.72 0.735 0.72 0.735 0.765 1.335 0.765 1.335 0.715 1.575 0.715 1.575 0.765 2.175 0.765 2.175 0.715 2.415 0.715 2.415 0.765 3.015 0.765 3.015 0.715 3.255 0.715 3.255 0.765 3.855 0.765 3.855 0.715 4.095 0.715 4.095 0.765 4.695 0.765 4.695 0.715 4.935 0.715 4.935 0.765 5.535 0.765 5.535 0.715 5.775 0.715 ;
  END
END NAND4X8

MACRO NOR4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX2 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.94 0.855 1.105 ;
        RECT 0.495 0.985 0.615 1.265 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 1.34 1.095 1.46 ;
        RECT 0.975 1.22 1.095 1.46 ;
        RECT 0.595 1.52 0.855 1.67 ;
        RECT 0.735 1.34 0.855 1.67 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.045 3.835 1.435 ;
        RECT 3.715 1.035 3.835 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 1.225 4.735 1.35 ;
        RECT 4.075 1.225 4.44 1.38 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.855 0.885 5.15 1.145 ;
        RECT 4.855 0.71 4.975 1.62 ;
        RECT 4.835 1.5 4.955 2.01 ;
        RECT 2.995 0.76 4.975 0.88 ;
        RECT 4.63 0.71 4.975 0.88 ;
        RECT 4.675 0.59 4.795 0.88 ;
        RECT 3.835 0.59 3.955 0.88 ;
        RECT 2.095 0.7 3.115 0.77 ;
        RECT 2.995 0.59 3.115 0.88 ;
        RECT 2.215 0.76 4.975 0.82 ;
        RECT 2.095 0.65 2.335 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 5.095 -0.18 5.215 0.64 ;
        RECT 4.255 -0.18 4.375 0.64 ;
        RECT 3.415 -0.18 3.535 0.64 ;
        RECT 2.515 0.46 2.755 0.58 ;
        RECT 2.515 -0.18 2.635 0.58 ;
        RECT 1.735 -0.18 1.855 0.64 ;
        RECT 0.715 -0.18 0.835 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 1.925 1.66 2.045 2.79 ;
        RECT 0.715 1.79 0.835 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.375 2.15 5.33 2.15 5.33 2.25 3.575 2.25 3.575 1.795 3.695 1.795 3.695 2.13 4.415 2.13 4.415 1.5 4.535 1.5 4.535 2.13 5.21 2.13 5.21 2.03 5.255 2.03 5.255 1.5 5.375 1.5 ;
      POLYGON 4.115 2.01 3.995 2.01 3.995 1.675 2.885 1.675 2.885 2.01 2.765 2.01 2.765 1.555 3.995 1.555 3.995 1.5 4.115 1.5 ;
      POLYGON 3.305 2.21 3.26 2.21 3.26 2.25 2.345 2.25 2.345 1.54 1.67 1.54 1.67 2.09 1.625 2.09 1.625 2.21 1.505 2.21 1.505 1.97 1.55 1.97 1.55 1.42 2.465 1.42 2.465 2.13 3.14 2.13 3.14 2.09 3.185 2.09 3.185 1.795 3.305 1.795 ;
      POLYGON 2.915 1.12 2.675 1.12 2.675 1.06 1.855 1.06 1.855 0.88 1.495 0.88 1.495 0.48 1.075 0.48 1.075 0.82 0.355 0.82 0.355 1.82 0.235 1.82 0.235 0.6 0.355 0.6 0.355 0.7 0.955 0.7 0.955 0.36 1.615 0.36 1.615 0.76 1.975 0.76 1.975 0.94 2.795 0.94 2.795 1 2.915 1 ;
      POLYGON 2.075 1.3 1.335 1.3 1.335 1.7 1.315 1.7 1.315 1.82 1.195 1.82 1.195 1.58 1.215 1.58 1.215 0.84 1.195 0.84 1.195 0.6 1.315 0.6 1.315 0.72 1.335 0.72 1.335 1.18 2.075 1.18 ;
  END
END NOR4BBX2

MACRO DFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX1 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 1.34 2.14 1.46 ;
        RECT 2.02 1.22 2.14 1.46 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.84 1.34 1.96 1.725 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.08 1.09 7.2 1.33 ;
        RECT 6.74 1.175 7.2 1.295 ;
        RECT 6.74 1.175 6.89 1.435 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.41 1.01 7.56 1.25 ;
        RECT 7.32 0.885 7.495 1.145 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.38 1.3 1.5 2.21 ;
        RECT 1.38 0.62 1.5 0.86 ;
        RECT 1.36 0.74 1.48 1.42 ;
        RECT 1.23 0.885 1.48 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 6.96 -0.18 7.08 0.91 ;
        RECT 4.83 -0.18 5.07 0.32 ;
        RECT 3.23 -0.18 3.35 0.9 ;
        RECT 1.8 -0.18 1.92 0.73 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.8 1.81 7.92 2.79 ;
        RECT 6.9 2.23 7.02 2.79 ;
        RECT 4.83 2.16 5.07 2.28 ;
        RECT 4.83 2.16 4.95 2.79 ;
        RECT 3.11 2.16 3.35 2.28 ;
        RECT 3.11 2.16 3.23 2.79 ;
        RECT 1.8 1.845 1.92 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.8 1.49 7.5 1.49 7.5 2.11 6.055 2.11 6.055 1.98 6.03 1.98 6.03 1.51 6.19 1.51 6.19 0.9 6.13 0.9 6.13 0.66 6.25 0.66 6.25 0.78 6.31 0.78 6.31 1.63 6.15 1.63 6.15 1.86 6.175 1.86 6.175 1.99 7.38 1.99 7.38 1.37 7.68 1.37 7.68 0.67 7.8 0.67 ;
      POLYGON 6.66 0.91 6.62 0.91 6.62 1.87 6.36 1.87 6.36 1.75 6.5 1.75 6.5 0.79 6.54 0.79 6.54 0.67 6.43 0.67 6.43 0.54 6.01 0.54 6.01 1.27 6.07 1.27 6.07 1.39 5.83 1.39 5.83 1.27 5.89 1.27 5.89 0.54 5.31 0.54 5.31 0.56 4.23 0.56 4.23 1 4.37 1 4.37 1.24 4.23 1.24 4.23 1.4 3.83 1.4 3.83 1.52 3.71 1.52 3.71 1.28 4.11 1.28 4.11 0.44 5.19 0.44 5.19 0.42 5.37 0.42 5.37 0.38 5.61 0.38 5.61 0.42 6.55 0.42 6.55 0.55 6.66 0.55 ;
      POLYGON 5.77 0.84 5.71 0.84 5.71 1.62 5.73 1.62 5.73 1.86 5.61 1.86 5.61 1.74 5.59 1.74 5.59 1.48 4.73 1.48 4.73 1.36 5.59 1.36 5.59 0.84 5.53 0.84 5.53 0.72 5.77 0.72 ;
      POLYGON 5.63 2.24 5.195 2.24 5.195 2.04 4.255 2.04 4.255 2.24 4.015 2.24 4.015 2.04 2.28 2.04 2.28 0.68 2.4 0.68 2.4 1.92 5.315 1.92 5.315 2.12 5.63 2.12 ;
      POLYGON 5.27 1.16 4.61 1.16 4.61 1.8 4.35 1.8 4.35 1.68 4.49 1.68 4.49 0.84 4.35 0.84 4.35 0.72 4.61 0.72 4.61 1.04 5.27 1.04 ;
      POLYGON 4.05 1.8 3.81 1.8 3.81 1.76 3.47 1.76 3.47 1.4 2.95 1.4 2.95 1.52 2.83 1.52 2.83 1.28 3.47 1.28 3.47 1.04 3.87 1.04 3.87 0.66 3.99 0.66 3.99 1.16 3.59 1.16 3.59 1.64 3.93 1.64 3.93 1.68 4.05 1.68 ;
      POLYGON 3.35 1.16 2.71 1.16 2.71 1.68 2.87 1.68 2.87 1.8 2.59 1.8 2.59 0.78 2.67 0.78 2.67 0.66 2.57 0.66 2.57 0.56 2.16 0.56 2.16 1.1 1.84 1.1 1.84 1.18 1.6 1.18 1.6 0.98 2.04 0.98 2.04 0.44 2.69 0.44 2.69 0.54 2.79 0.54 2.79 0.9 2.71 0.9 2.71 1.04 3.35 1.04 ;
      POLYGON 1.11 1.08 1.095 1.08 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.96 0.99 0.96 0.99 0.68 1.11 0.68 ;
  END
END DFFTRX1

MACRO TLATXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATXL 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.03 0.85 1.435 ;
        RECT 0.73 1.015 0.85 1.435 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.14 3.41 1.59 ;
        RECT 3.26 1.14 3.38 1.615 ;
    END
  END G
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.01 0.54 4.13 0.78 ;
        RECT 3.84 1.465 4.08 1.735 ;
        RECT 3.96 0.66 4.08 1.735 ;
        RECT 3.81 1.615 3.93 1.855 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.24 0.62 5.36 1.175 ;
        RECT 5.04 1.055 5.36 1.175 ;
        RECT 5.04 1.055 5.16 1.72 ;
        RECT 5 1.175 5.16 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.82 -0.18 4.94 0.86 ;
        RECT 3.59 -0.18 3.71 0.78 ;
        RECT 2.3 -0.18 2.42 0.395 ;
        RECT 0.615 -0.18 0.735 0.395 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.62 1.6 4.74 2.79 ;
        RECT 3.39 1.735 3.51 2.79 ;
        RECT 1.93 2.215 2.17 2.79 ;
        RECT 0.59 1.795 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.88 1.34 4.5 1.34 4.5 1.6 4.32 1.6 4.32 1.72 4.2 1.72 4.2 1.48 4.38 1.48 4.38 1.1 4.4 1.1 4.4 0.62 4.52 0.62 4.52 1.22 4.88 1.22 ;
      POLYGON 3.84 1.06 3.6 1.06 3.6 1.02 2.9 1.02 2.9 1.515 2.65 1.515 2.65 1.855 2.41 1.855 2.41 1.735 2.53 1.735 2.53 1.515 1.93 1.515 1.93 1.395 2.78 1.395 2.78 0.675 2.9 0.675 2.9 0.9 3.84 0.9 ;
      POLYGON 3.29 0.78 3.17 0.78 3.17 0.555 2.66 0.555 2.66 0.635 2.01 0.635 2.01 0.615 1.43 0.615 1.43 1.475 1.21 1.475 1.21 1.595 1.11 1.595 1.11 2.075 1.52 2.075 1.52 1.975 2.97 1.975 2.97 1.735 3.09 1.735 3.09 2.095 1.64 2.095 1.64 2.195 0.99 2.195 0.99 1.675 0.41 1.675 0.41 1.335 0.53 1.335 0.53 1.555 0.99 1.555 0.99 1.355 1.31 1.355 1.31 0.495 1.71 0.495 1.71 0.395 1.95 0.395 1.95 0.495 2.13 0.495 2.13 0.515 2.54 0.515 2.54 0.435 3.29 0.435 ;
      POLYGON 2.49 1.275 1.67 1.275 1.67 1.835 1.35 1.835 1.35 1.955 1.23 1.955 1.23 1.715 1.55 1.715 1.55 0.735 1.79 0.735 1.79 0.855 1.67 0.855 1.67 1.155 2.49 1.155 ;
      POLYGON 1.19 1.235 1.07 1.235 1.07 0.895 0.29 0.895 0.29 1.915 0.17 1.915 0.17 0.915 0.135 0.915 0.135 0.675 0.255 0.675 0.255 0.775 1.19 0.775 ;
  END
END TLATXL

MACRO AO22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X4 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.815 0.82 1.235 ;
        RECT 0.7 0.795 0.82 1.235 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.055 0.905 1.175 1.235 ;
        RECT 0.94 0.885 1.09 1.215 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.76 0.51 1.21 ;
        RECT 0.38 0.76 0.5 1.235 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.23 2.015 1.38 ;
        RECT 1.535 1.17 1.875 1.29 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 1.175 3.7 1.435 ;
        RECT 2.545 1.32 3.525 1.44 ;
        RECT 3.405 0.69 3.525 1.44 ;
        RECT 3.385 1.32 3.505 2.21 ;
        RECT 2.155 0.69 3.525 0.81 ;
        RECT 2.995 0.65 3.235 0.81 ;
        RECT 2.545 1.32 2.665 2.21 ;
        RECT 2.035 0.65 2.275 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.475 0.45 3.715 0.57 ;
        RECT 3.475 -0.18 3.595 0.57 ;
        RECT 2.515 0.45 2.755 0.57 ;
        RECT 2.515 -0.18 2.635 0.57 ;
        RECT 1.675 -0.18 1.795 0.64 ;
        RECT 0.22 -0.18 0.34 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 3.805 1.56 3.925 2.79 ;
        RECT 2.965 1.56 3.085 2.79 ;
        RECT 2.065 2.23 2.185 2.79 ;
        RECT 0.555 1.595 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.285 1.09 3.045 1.09 3.045 1.05 2.535 1.05 2.535 1.11 2.295 1.11 2.295 1.05 1.415 1.05 1.415 1.41 1.515 1.41 1.515 2.01 1.395 2.01 1.395 1.53 1.295 1.53 1.295 0.675 0.915 0.675 0.915 0.555 1.415 0.555 1.415 0.93 3.165 0.93 3.165 0.97 3.285 0.97 ;
      POLYGON 1.935 2.25 0.975 2.25 0.975 1.475 0.255 1.475 0.255 2.08 0.135 2.08 0.135 1.355 1.095 1.355 1.095 2.13 1.815 2.13 1.815 1.5 1.935 1.5 ;
  END
END AO22X4

MACRO NAND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X6 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.075 1.17 7.735 1.29 ;
        RECT 6.975 1.23 7.235 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.29 1.175 5.595 1.33 ;
        RECT 5.475 1.09 5.595 1.33 ;
        RECT 5.29 1.175 5.44 1.435 ;
        RECT 5.095 1.15 5.335 1.27 ;
        RECT 5.215 1.175 5.595 1.295 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.295 1.17 3.535 1.29 ;
        RECT 2.97 1.175 3.415 1.295 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 2.995 1.11 3.115 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.175 1.38 1.435 ;
        RECT 1.255 1.11 1.375 1.435 ;
        RECT 0.955 1.175 1.38 1.295 ;
        RECT 0.835 1.17 1.075 1.29 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.9712 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.995 0.93 8.855 1.05 ;
        RECT 8.735 0.4 8.855 1.05 ;
        RECT 8.255 1.43 8.375 2.21 ;
        RECT 0.695 1.555 8.375 1.675 ;
        RECT 7.9 1.175 8.05 1.435 ;
        RECT 7.9 0.93 8.02 1.675 ;
        RECT 7.835 0.6 7.955 1.05 ;
        RECT 7.415 1.43 7.535 2.21 ;
        RECT 6.995 0.6 7.115 1.05 ;
        RECT 6.575 1.43 6.695 2.21 ;
        RECT 5.735 1.43 5.855 2.21 ;
        RECT 4.895 1.43 5.015 2.21 ;
        RECT 4.055 1.43 4.175 2.21 ;
        RECT 3.215 1.555 3.335 2.21 ;
        RECT 2.375 1.43 2.495 2.21 ;
        RECT 1.535 1.43 1.655 2.21 ;
        RECT 0.695 1.43 0.815 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 1.875 -0.18 1.995 0.75 ;
        RECT 1.035 -0.18 1.155 0.75 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.675 1.43 8.795 2.79 ;
        RECT 7.835 1.795 7.955 2.79 ;
        RECT 6.995 1.795 7.115 2.79 ;
        RECT 6.155 1.795 6.275 2.79 ;
        RECT 5.315 1.795 5.435 2.79 ;
        RECT 4.475 1.795 4.595 2.79 ;
        RECT 3.635 1.795 3.755 2.79 ;
        RECT 2.795 1.795 2.915 2.79 ;
        RECT 1.955 1.795 2.075 2.79 ;
        RECT 1.115 1.795 1.235 2.79 ;
        RECT 0.275 1.43 0.395 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.435 0.81 8.315 0.81 8.315 0.48 7.535 0.48 7.535 0.81 7.415 0.81 7.415 0.48 6.695 0.48 6.695 0.92 6.575 0.92 6.575 0.48 5.855 0.48 5.855 0.73 5.735 0.73 5.735 0.48 4.955 0.48 4.955 0.73 4.835 0.73 4.835 0.36 8.435 0.36 ;
      POLYGON 6.275 0.97 4.415 0.97 4.415 0.48 3.675 0.48 3.675 0.75 3.555 0.75 3.555 0.48 2.835 0.48 2.835 0.75 2.715 0.75 2.715 0.36 4.535 0.36 4.535 0.85 5.315 0.85 5.315 0.6 5.435 0.6 5.435 0.85 6.155 0.85 6.155 0.6 6.275 0.6 ;
      POLYGON 4.115 0.99 0.555 0.99 0.555 0.4 0.675 0.4 0.675 0.87 1.455 0.87 1.455 0.4 1.575 0.4 1.575 0.87 2.295 0.87 2.295 0.4 2.415 0.4 2.415 0.87 3.135 0.87 3.135 0.6 3.255 0.6 3.255 0.87 3.995 0.87 3.995 0.6 4.115 0.6 ;
  END
END NAND4X6

MACRO SDFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX2 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.275 0.36 6.515 0.48 ;
        RECT 5.695 0.85 6.415 0.97 ;
        RECT 6.295 0.36 6.415 0.97 ;
        RECT 5.695 0.38 5.815 0.97 ;
        RECT 4.365 0.36 5.81 0.48 ;
        RECT 5.69 0.38 5.815 0.5 ;
        RECT 4.365 1.23 4.625 1.38 ;
        RECT 4.365 0.36 4.485 1.38 ;
        RECT 3.685 1.24 4.625 1.36 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.145 0.845 9.465 1.01 ;
        RECT 9.005 0.89 9.265 1.09 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.585 0.775 9.825 0.98 ;
        RECT 9.64 0.76 9.79 1.155 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.785 1.26 11.295 1.385 ;
        RECT 11.035 1.23 11.295 1.385 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.185 0.925 11.225 1.045 ;
        RECT 10.745 0.925 11.005 1.09 ;
        RECT 10.445 0.76 10.565 1.045 ;
        RECT 10.065 1.515 10.305 1.635 ;
        RECT 10.185 0.925 10.305 1.635 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.59 0.675 2.21 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.195 0.68 2.315 1.99 ;
        RECT 2.1 1.175 2.315 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.925 -0.18 11.045 0.64 ;
        RECT 9.645 -0.18 9.765 0.64 ;
        RECT 7.355 -0.18 7.475 0.58 ;
        RECT 5.935 0.61 6.175 0.73 ;
        RECT 6.035 -0.18 6.155 0.73 ;
        RECT 3.525 0.66 3.765 0.78 ;
        RECT 3.525 -0.18 3.645 0.78 ;
        RECT 2.615 -0.18 2.735 0.78 ;
        RECT 1.775 -0.18 1.895 0.73 ;
        RECT 1.035 -0.18 1.155 0.53 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 10.925 1.935 11.045 2.79 ;
        RECT 9.585 1.995 9.825 2.115 ;
        RECT 9.585 1.995 9.705 2.79 ;
        RECT 7.455 1.66 7.575 2.79 ;
        RECT 6.435 2.29 6.675 2.79 ;
        RECT 4.185 2.05 4.425 2.17 ;
        RECT 4.185 2.05 4.305 2.79 ;
        RECT 3.345 1.97 3.465 2.79 ;
        RECT 2.675 2.14 2.795 2.79 ;
        RECT 1.715 1.98 1.835 2.79 ;
        RECT 0.975 1.73 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.535 1.745 11.465 1.745 11.465 2.055 11.345 2.055 11.345 1.625 10.545 1.625 10.545 1.375 10.425 1.375 10.425 1.255 10.665 1.255 10.665 1.505 11.415 1.505 11.415 1.11 11.345 1.11 11.345 0.4 11.465 0.4 11.465 0.99 11.535 0.99 ;
      POLYGON 10.405 0.64 10.065 0.64 10.065 1.395 9.945 1.395 9.945 1.755 10.405 1.755 10.405 2.055 10.285 2.055 10.285 1.875 8.755 1.875 8.755 1.76 8.635 1.76 8.635 1.64 8.755 1.64 8.755 0.72 8.695 0.72 8.695 0.6 8.935 0.6 8.935 0.72 8.875 0.72 8.875 1.755 9.825 1.755 9.825 1.275 9.945 1.275 9.945 0.52 10.285 0.52 10.285 0.4 10.405 0.4 ;
      POLYGON 9.405 2.115 8.395 2.115 8.395 1.99 8.175 1.99 8.175 2.15 7.935 2.15 7.935 1.99 7.745 1.99 7.745 1.54 7.335 1.54 7.335 2.11 6.805 2.11 6.805 2.17 6.115 2.17 6.115 2.05 6.685 2.05 6.685 1.99 7.215 1.99 7.215 1.42 7.865 1.42 7.865 1.87 8.395 1.87 8.395 1.4 8.455 1.4 8.455 0.36 9.265 0.36 9.265 0.64 9.145 0.64 9.145 0.48 8.575 0.48 8.575 1.52 8.515 1.52 8.515 1.995 9.405 1.995 ;
      POLYGON 8.335 1.28 8.275 1.28 8.275 1.75 8.155 1.75 8.155 1.3 7.175 1.3 7.175 1.18 8.155 1.18 8.155 1.16 8.215 1.16 8.215 0.72 8.095 0.72 8.095 0.6 8.335 0.6 ;
      POLYGON 8.095 1.04 7.855 1.04 7.855 0.82 7.115 0.82 7.115 0.5 6.755 0.5 6.755 0.72 6.655 0.72 6.655 1.21 6.075 1.21 6.075 1.57 6.195 1.57 6.195 1.69 5.955 1.69 5.955 1.21 5.225 1.21 5.225 1.03 5.455 1.03 5.455 0.62 5.575 0.62 5.575 1.09 6.535 1.09 6.535 0.6 6.635 0.6 6.635 0.38 7.235 0.38 7.235 0.7 7.975 0.7 7.975 0.92 8.095 0.92 ;
      POLYGON 7.735 1.06 6.995 1.06 6.995 1.51 7.095 1.51 7.095 1.87 6.565 1.87 6.565 1.93 5.625 1.93 5.625 1.45 4.985 1.45 4.985 0.72 5.025 0.72 5.025 0.6 5.145 0.6 5.145 0.84 5.105 0.84 5.105 1.33 5.745 1.33 5.745 1.81 6.445 1.81 6.445 1.75 6.975 1.75 6.975 1.63 6.875 1.63 6.875 0.62 6.995 0.62 6.995 0.94 7.735 0.94 ;
      POLYGON 5.325 1.87 5.205 1.87 5.205 1.69 3.445 1.69 3.445 1.38 3.275 1.38 3.275 1.14 3.395 1.14 3.395 1.26 3.565 1.26 3.565 1.57 4.745 1.57 4.745 1.11 4.605 1.11 4.605 0.6 4.725 0.6 4.725 0.99 4.865 0.99 4.865 1.57 5.325 1.57 ;
      POLYGON 4.965 1.93 3.945 1.93 3.945 2.03 3.705 2.03 3.705 1.91 3.825 1.91 3.825 1.81 4.965 1.81 ;
      POLYGON 4.245 1.12 4.005 1.12 4.005 1.02 3.155 1.02 3.155 1.82 3.035 1.82 3.035 1.02 2.595 1.02 2.595 1.24 2.475 1.24 2.475 0.9 3.035 0.9 3.035 0.64 3.155 0.64 3.155 0.9 4.125 0.9 4.125 1 4.245 1 ;
      POLYGON 1.415 1.05 1.405 1.05 1.405 1.58 1.285 1.58 1.285 1.17 0.795 1.17 0.795 1.05 1.285 1.05 1.285 0.93 1.295 0.93 1.295 0.68 1.415 0.68 ;
  END
END SDFFSX2

MACRO MX3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X2 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.23 1.265 1.39 ;
        RECT 1.145 1.13 1.265 1.39 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.71 0.76 2.83 1.43 ;
        RECT 2.68 0.76 2.83 1.16 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.885 3.315 1.06 ;
        RECT 3.195 0.82 3.315 1.06 ;
        RECT 2.97 0.885 3.12 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.42 1.085 4.57 1.46 ;
        RECT 4.295 1.11 4.57 1.3 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.71 1.465 4.86 1.725 ;
        RECT 4.71 1.46 4.83 1.725 ;
        RECT 4.015 1.58 4.86 1.7 ;
        RECT 4.015 1.46 4.135 1.7 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 1.35 0.765 2.16 ;
        RECT 0.485 0.65 0.765 0.77 ;
        RECT 0.645 0.53 0.765 0.77 ;
        RECT 0.485 1.35 0.765 1.47 ;
        RECT 0.305 1.23 0.605 1.38 ;
        RECT 0.485 0.65 0.605 1.47 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 4.415 -0.18 4.535 0.64 ;
        RECT 3.135 -0.18 3.255 0.64 ;
        RECT 1.005 0.48 1.245 0.6 ;
        RECT 1.005 -0.18 1.125 0.6 ;
        RECT 0.225 -0.18 0.345 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.515 1.94 4.635 2.79 ;
        RECT 3.195 1.94 3.315 2.79 ;
        RECT 1.065 1.51 1.185 2.79 ;
        RECT 0.225 1.51 0.345 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.1 1.965 5.055 1.965 5.055 2.085 4.935 2.085 4.935 1.845 4.98 1.845 4.98 0.965 4.055 0.965 4.055 1 3.895 1 3.895 1.46 3.795 1.46 3.795 1.58 3.675 1.58 3.675 1.34 3.775 1.34 3.775 0.845 3.935 0.845 3.935 0.76 4.055 0.76 4.055 0.845 4.98 0.845 4.98 0.64 4.835 0.64 4.835 0.4 4.955 0.4 4.955 0.52 5.1 0.52 ;
      POLYGON 3.955 2.06 3.835 2.06 3.835 1.94 3.775 1.94 3.775 1.82 2.405 1.82 2.405 1.69 2.185 1.69 2.185 1.57 2.405 1.57 2.405 0.79 2.265 0.79 2.265 0.67 2.525 0.67 2.525 1.7 3.435 1.7 3.435 1.1 3.535 1.1 3.535 0.52 3.775 0.52 3.775 0.4 3.895 0.4 3.895 0.64 3.655 0.64 3.655 1.22 3.555 1.22 3.555 1.7 3.895 1.7 3.895 1.82 3.955 1.82 ;
      POLYGON 2.955 2.06 1.945 2.06 1.945 1.29 1.745 1.29 1.745 1.41 1.625 1.41 1.625 1.17 2.165 1.17 2.165 1.03 2.025 1.03 2.025 0.43 2.715 0.43 2.715 0.4 2.835 0.4 2.835 0.64 2.715 0.64 2.715 0.55 2.145 0.55 2.145 0.91 2.285 0.91 2.285 1.45 2.065 1.45 2.065 1.94 2.955 1.94 ;
      POLYGON 1.905 1.01 1.505 1.01 1.505 1.53 1.825 1.53 1.825 1.77 1.705 1.77 1.705 1.65 1.385 1.65 1.385 1.01 0.965 1.01 0.965 1.11 0.725 1.11 0.725 0.89 1.785 0.89 1.785 0.61 1.905 0.61 ;
  END
END MX3X2

MACRO NOR4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX2 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.175 4.12 1.385 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 1.23 3.525 1.4 ;
        RECT 3.195 1.1 3.355 1.38 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.385 1.29 2.885 1.41 ;
        RECT 2.625 1.18 2.885 1.41 ;
        RECT 2.385 1 2.505 1.41 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.395 1.295 ;
        RECT 0.275 1.055 0.395 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.195 1.53 4.315 2.01 ;
        RECT 2.145 1.53 4.315 1.65 ;
        RECT 1.305 0.76 3.945 0.88 ;
        RECT 3.825 0.59 3.945 0.88 ;
        RECT 2.985 0.59 3.105 0.88 ;
        RECT 2.145 0.59 2.265 1.65 ;
        RECT 2.1 1.175 2.265 1.435 ;
        RECT 1.305 0.59 1.425 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.245 -0.18 4.365 0.64 ;
        RECT 3.405 -0.18 3.525 0.64 ;
        RECT 2.565 -0.18 2.685 0.64 ;
        RECT 1.725 -0.18 1.845 0.64 ;
        RECT 0.825 -0.18 0.945 0.53 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 1.225 2.01 1.465 2.15 ;
        RECT 1.225 2.01 1.345 2.79 ;
        RECT 0.135 1.555 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.735 2.25 3.775 2.25 3.775 1.89 3.055 1.89 3.055 2.01 2.935 2.01 2.935 1.77 3.895 1.77 3.895 2.13 4.615 2.13 4.615 1.56 4.735 1.56 ;
      POLYGON 3.535 2.15 3.415 2.15 3.415 2.25 2.185 2.25 2.185 2.15 2.065 2.15 2.065 2.01 2.305 2.01 2.305 2.13 3.295 2.13 3.295 2.01 3.535 2.01 ;
      POLYGON 2.665 2.01 2.545 2.01 2.545 1.89 1.825 1.89 1.825 2.21 1.705 2.21 1.705 1.89 0.985 1.89 0.985 2.21 0.865 2.21 0.865 1.77 1.705 1.77 1.705 1.56 1.825 1.56 1.825 1.77 2.665 1.77 ;
      POLYGON 1.225 1.19 0.675 1.19 0.675 1.675 0.555 1.675 0.555 0.68 0.675 0.68 0.675 1.07 1.225 1.07 ;
  END
END NOR4BX2

MACRO OAI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222XL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.14 1.96 1.61 ;
    END
  END B0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.14 2.83 1.61 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.14 0.885 1.47 ;
        RECT 0.65 1.14 0.8 1.475 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.16 2.375 1.28 ;
        RECT 2.255 1.025 2.375 1.28 ;
        RECT 2.1 1.16 2.25 1.435 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.14 0.51 1.515 ;
        RECT 0.39 0.96 0.51 1.515 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 1.15 1.67 1.61 ;
        RECT 1.515 1.14 1.635 1.61 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4116 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.73 3.07 1.85 ;
        RECT 2.95 0.9 3.07 1.85 ;
        RECT 2.635 0.9 3.07 1.02 ;
        RECT 2.735 1.73 2.855 2.09 ;
        RECT 2.635 0.72 2.755 1.02 ;
        RECT 2.68 1.73 2.855 2.015 ;
        RECT 2.515 0.6 2.635 0.84 ;
        RECT 1.255 1.73 1.375 2.09 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 0.985 -0.18 1.105 0.45 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.095 1.97 2.215 2.79 ;
        RECT 0.285 1.97 0.405 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.115 0.78 2.875 0.78 2.875 0.48 2.215 0.48 2.215 0.84 2.095 0.84 2.095 0.48 1.435 0.48 1.435 0.78 1.195 0.78 1.195 0.66 1.315 0.66 1.315 0.36 2.995 0.36 2.995 0.66 3.115 0.66 ;
      POLYGON 1.795 1.02 0.63 1.02 0.63 0.84 0.445 0.84 0.445 0.72 0.75 0.72 0.75 0.9 1.675 0.9 1.675 0.6 1.795 0.6 ;
  END
END OAI222XL

MACRO AOI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X4 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.275 1.02 3.515 1.14 ;
        RECT 0.515 0.99 3.395 1.11 ;
        RECT 1.995 0.99 2.235 1.14 ;
        RECT 0.595 0.94 0.855 1.11 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.625 0.99 10.505 1.11 ;
        RECT 10.165 0.94 10.425 1.11 ;
        RECT 8.785 0.99 9.025 1.14 ;
        RECT 7.505 1.02 7.745 1.14 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.005 1.02 7.245 1.14 ;
        RECT 4.365 0.99 7.125 1.11 ;
        RECT 5.455 0.99 5.695 1.14 ;
        RECT 4.365 1.23 4.625 1.38 ;
        RECT 4.365 0.99 4.485 1.38 ;
        RECT 4.165 1.02 4.485 1.14 ;
    END
  END B0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.145 1.26 9.665 1.38 ;
        RECT 9.295 1.23 9.555 1.38 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.355 1.26 2.875 1.38 ;
        RECT 1.465 1.23 1.725 1.38 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.905 1.26 6.405 1.38 ;
        RECT 5.815 1.23 6.075 1.38 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.6576 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.265 1.5 10.385 2.01 ;
        RECT 3.925 1.5 10.385 1.62 ;
        RECT 9.425 1.5 9.545 2.01 ;
        RECT 9.265 0.68 9.505 0.8 ;
        RECT 1.635 0.73 9.385 0.85 ;
        RECT 8.585 1.5 8.705 2.01 ;
        RECT 7.985 0.68 8.225 0.85 ;
        RECT 7.745 1.5 7.865 2.01 ;
        RECT 6.425 0.68 6.665 0.85 ;
        RECT 4.645 0.68 4.885 0.85 ;
        RECT 3.925 0.73 4.045 1.62 ;
        RECT 3.785 1.23 4.045 1.38 ;
        RECT 2.795 0.68 3.035 0.85 ;
        RECT 1.515 0.68 1.755 0.8 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 9.965 -0.18 10.085 0.67 ;
        RECT 8.625 0.49 8.865 0.61 ;
        RECT 8.625 -0.18 8.745 0.61 ;
        RECT 7.265 0.49 7.505 0.61 ;
        RECT 7.265 -0.18 7.385 0.61 ;
        RECT 5.385 0.49 5.625 0.61 ;
        RECT 5.385 -0.18 5.505 0.61 ;
        RECT 3.905 0.49 4.145 0.61 ;
        RECT 3.905 -0.18 4.025 0.61 ;
        RECT 2.155 0.49 2.395 0.61 ;
        RECT 2.155 -0.18 2.275 0.61 ;
        RECT 0.935 -0.18 1.055 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 3.515 1.98 3.755 2.15 ;
        RECT 3.515 1.98 3.635 2.79 ;
        RECT 2.675 1.98 2.915 2.15 ;
        RECT 2.675 1.98 2.795 2.79 ;
        RECT 1.835 1.98 2.075 2.15 ;
        RECT 1.835 1.98 1.955 2.79 ;
        RECT 0.995 1.98 1.235 2.15 ;
        RECT 0.995 1.98 1.115 2.79 ;
        RECT 0.215 1.56 0.335 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.805 2.25 4.025 2.25 4.025 2.15 3.905 2.15 3.905 1.98 4.145 1.98 4.145 2.13 4.745 2.13 4.745 1.98 4.985 1.98 4.985 2.13 5.585 2.13 5.585 1.98 5.825 1.98 5.825 2.13 6.425 2.13 6.425 1.98 6.665 1.98 6.665 2.13 7.325 2.13 7.325 1.74 7.445 1.74 7.445 2.13 8.165 2.13 8.165 1.74 8.285 1.74 8.285 2.13 9.005 2.13 9.005 1.74 9.125 1.74 9.125 2.13 9.845 2.13 9.845 1.74 9.965 1.74 9.965 2.13 10.685 2.13 10.685 1.56 10.805 1.56 ;
      POLYGON 7.025 2.01 6.905 2.01 6.905 1.86 6.185 1.86 6.185 2.01 6.065 2.01 6.065 1.86 5.345 1.86 5.345 2.01 5.225 2.01 5.225 1.86 4.505 1.86 4.505 2.01 4.385 2.01 4.385 1.86 3.275 1.86 3.275 2.21 3.155 2.21 3.155 1.86 2.435 1.86 2.435 2.21 2.315 2.21 2.315 1.86 1.595 1.86 1.595 2.21 1.475 2.21 1.475 1.86 0.755 1.86 0.755 2.21 0.635 2.21 0.635 1.56 0.755 1.56 0.755 1.74 1.475 1.74 1.475 1.56 1.595 1.56 1.595 1.74 2.315 1.74 2.315 1.56 2.435 1.56 2.435 1.74 3.155 1.74 3.155 1.56 3.275 1.56 3.275 1.74 7.025 1.74 ;
  END
END AOI222X4

MACRO CLKINVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX6 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.15 1.4 1.27 ;
        RECT 0.885 1.15 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.32 1.43 2.44 2.21 ;
        RECT 0.58 0.91 2.44 1.03 ;
        RECT 2.32 0.4 2.44 1.03 ;
        RECT 0.64 1.5 2.44 1.62 ;
        RECT 1.52 1.175 1.67 1.62 ;
        RECT 1.52 0.91 1.64 1.62 ;
        RECT 1.48 1.43 1.6 2.21 ;
        RECT 1.48 0.4 1.6 1.03 ;
        RECT 0.64 1.43 0.76 2.21 ;
        RECT 0.58 0.4 0.7 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.9 -0.18 2.02 0.79 ;
        RECT 1.06 -0.18 1.18 0.79 ;
        RECT 0.16 -0.18 0.28 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.9 1.74 2.02 2.79 ;
        RECT 1.06 1.74 1.18 2.79 ;
        RECT 0.22 1.43 0.34 2.79 ;
    END
  END VDD
END CLKINVX6

MACRO NOR4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX4 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.645 1.26 7.565 1.38 ;
        RECT 6.645 1.23 6.945 1.38 ;
        RECT 6.645 1 6.765 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 1.26 5.885 1.38 ;
        RECT 4.965 1.23 5.565 1.35 ;
        RECT 4.965 1 5.085 1.35 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 1.23 3.785 1.35 ;
        RECT 3.205 1.23 3.465 1.38 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 1 0.395 1.24 ;
        RECT 0.07 1 0.395 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.645 1.5 7.765 2.01 ;
        RECT 2.965 1.5 7.765 1.62 ;
        RECT 1.345 0.76 7.345 0.88 ;
        RECT 7.225 0.59 7.345 0.88 ;
        RECT 6.805 1.5 6.925 2.01 ;
        RECT 6.385 0.59 6.505 0.88 ;
        RECT 5.545 0.59 5.665 0.88 ;
        RECT 4.705 0.59 4.825 0.88 ;
        RECT 3.865 0.59 3.985 0.88 ;
        RECT 2.915 1.52 3.175 1.67 ;
        RECT 3.025 0.59 3.145 0.88 ;
        RECT 2.965 0.76 3.085 1.67 ;
        RECT 2.185 0.59 2.305 0.88 ;
        RECT 1.345 0.59 1.465 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.645 -0.18 7.765 0.64 ;
        RECT 6.805 -0.18 6.925 0.64 ;
        RECT 5.965 -0.18 6.085 0.64 ;
        RECT 5.125 -0.18 5.245 0.64 ;
        RECT 4.285 -0.18 4.405 0.64 ;
        RECT 3.445 -0.18 3.565 0.64 ;
        RECT 2.605 -0.18 2.725 0.64 ;
        RECT 1.765 -0.18 1.885 0.64 ;
        RECT 0.865 -0.18 0.985 0.53 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 2.125 2.03 2.365 2.15 ;
        RECT 2.125 2.03 2.245 2.79 ;
        RECT 1.285 2.03 1.525 2.15 ;
        RECT 1.285 2.03 1.405 2.79 ;
        RECT 0.135 1.36 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.185 2.25 6.385 2.25 6.385 1.86 5.725 1.86 5.725 2.01 5.485 2.01 5.485 1.86 4.885 1.86 4.885 2.01 4.645 2.01 4.645 1.74 6.505 1.74 6.505 2.13 7.225 2.13 7.225 1.74 7.345 1.74 7.345 2.13 8.065 2.13 8.065 1.56 8.185 1.56 ;
      POLYGON 6.145 2.15 6.025 2.15 6.025 2.25 3.085 2.25 3.085 2.15 2.965 2.15 2.965 2.03 3.205 2.03 3.205 2.13 3.805 2.13 3.805 2.03 4.045 2.03 4.045 2.13 5.065 2.13 5.065 1.98 5.305 1.98 5.305 2.13 5.905 2.13 5.905 1.98 6.145 1.98 ;
      POLYGON 4.465 2.01 4.225 2.01 4.225 1.91 3.625 1.91 3.625 2.01 3.385 2.01 3.385 1.91 2.725 1.91 2.725 2.21 2.605 2.21 2.605 1.91 1.885 1.91 1.885 2.21 1.765 2.21 1.765 1.91 1.045 1.91 1.045 2.21 0.925 2.21 0.925 1.79 1.765 1.79 1.765 1.56 1.885 1.56 1.885 1.79 2.605 1.79 2.605 1.56 2.725 1.56 2.725 1.79 3.385 1.79 3.385 1.74 3.625 1.74 3.625 1.79 4.225 1.79 4.225 1.74 4.465 1.74 ;
      POLYGON 2.105 1.32 0.675 1.32 0.675 1.64 0.555 1.64 0.555 0.68 0.675 0.68 0.675 1.2 2.105 1.2 ;
  END
END NOR4BX4

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.025 0.425 1.265 ;
        RECT 0.07 1.025 0.425 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.845 1.175 1.145 1.38 ;
        RECT 0.845 1.07 0.965 1.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.505 0.885 1.67 1.145 ;
        RECT 1.505 0.59 1.625 1.48 ;
        RECT 1.485 1.36 1.605 2.2 ;
        RECT 1.485 0.47 1.605 0.71 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 1.005 0.53 1.245 0.65 ;
        RECT 1.005 -0.18 1.125 0.65 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.065 1.55 1.185 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.385 1.24 1.265 1.24 1.265 0.95 0.705 0.95 0.705 1.505 0.545 1.505 0.545 1.73 0.305 1.73 0.305 1.61 0.425 1.61 0.425 1.385 0.585 1.385 0.585 0.66 0.705 0.66 0.705 0.83 1.385 0.83 ;
  END
END OR2X1

MACRO MX4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X4 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.455 1.57 3.695 1.69 ;
        RECT 3.435 0.74 3.675 0.86 ;
        RECT 3.455 0.74 3.575 1.69 ;
        RECT 2.68 1.315 3.575 1.435 ;
        RECT 2.535 1.175 2.83 1.315 ;
        RECT 2.495 1.57 2.8 1.69 ;
        RECT 2.68 1.175 2.8 1.69 ;
        RECT 2.535 0.68 2.655 1.315 ;
    END
  END Y
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.94 2.015 1.155 ;
        RECT 1.775 0.94 1.895 1.33 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 1.02 4.155 1.26 ;
        RECT 3.84 1.02 4.155 1.145 ;
        RECT 3.84 0.885 3.99 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 1.4 5.495 1.67 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 1.52 6.075 1.67 ;
        RECT 5.635 1.52 6.075 1.64 ;
        RECT 5.635 1.4 5.755 1.64 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.215 1.23 7.525 1.425 ;
        RECT 7.215 1.23 7.335 1.56 ;
    END
  END D
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2496 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.3867 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.9 1.175 8.05 1.435 ;
        RECT 7.645 1.1 8.02 1.22 ;
        RECT 7.645 0.99 7.765 1.34 ;
        RECT 6.795 0.99 7.765 1.11 ;
        RECT 6.795 0.99 6.915 1.24 ;
    END
  END S0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.235 0.74 7.475 0.86 ;
        RECT 7.235 -0.18 7.355 0.86 ;
        RECT 5.575 0.68 5.815 0.8 ;
        RECT 5.695 -0.18 5.815 0.8 ;
        RECT 4.035 -0.18 4.155 0.4 ;
        RECT 2.955 -0.18 3.195 0.32 ;
        RECT 1.995 -0.18 2.235 0.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.375 1.92 7.495 2.79 ;
        RECT 5.435 2.03 5.675 2.15 ;
        RECT 5.435 2.03 5.555 2.79 ;
        RECT 3.935 2.05 4.175 2.17 ;
        RECT 3.935 2.05 4.055 2.79 ;
        RECT 2.975 2.05 3.215 2.17 ;
        RECT 2.975 2.05 3.095 2.79 ;
        RECT 2.015 2.29 2.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.29 1.92 7.915 1.92 7.915 2.04 7.795 2.04 7.795 1.8 7.035 1.8 7.035 2.22 6.315 2.22 6.315 1.91 4.995 1.91 4.995 1.69 4.935 1.69 4.935 1.45 5.055 1.45 5.055 1.57 5.115 1.57 5.115 1.79 6.315 1.79 6.315 1.02 6.435 1.02 6.435 2.1 6.915 2.1 6.915 1.66 6.815 1.66 6.815 1.54 7.055 1.54 7.055 1.68 8.17 1.68 8.17 0.86 7.655 0.86 7.655 0.74 8.29 0.74 ;
      POLYGON 6.795 1.98 6.555 1.98 6.555 0.9 6.145 0.9 6.145 1.04 5.23 1.04 5.23 0.56 4.395 0.56 4.395 0.64 3.795 0.64 3.795 0.62 3 0.62 3 0.56 1.755 0.56 1.755 0.48 1.215 0.48 1.215 0.6 1.285 0.6 1.285 1.56 1.385 1.56 1.385 1.69 1.145 1.69 1.145 1.56 1.165 1.56 1.165 0.72 1.095 0.72 1.095 0.36 1.875 0.36 1.875 0.44 3.12 0.44 3.12 0.5 3.915 0.5 3.915 0.52 4.275 0.52 4.275 0.44 5.35 0.44 5.35 0.92 6.025 0.92 6.025 0.78 6.555 0.78 6.555 0.68 6.675 0.68 6.675 1.86 6.795 1.86 ;
      POLYGON 6.155 1.4 5.915 1.4 5.915 1.28 4.635 1.28 4.635 1.48 4.515 1.48 4.515 1.16 6.155 1.16 ;
      POLYGON 5.055 0.92 4.395 0.92 4.395 1.81 4.875 1.81 4.875 1.98 4.635 1.98 4.635 1.93 2.47 1.93 2.47 2.17 1.41 2.17 1.41 2.25 0.365 2.25 0.365 1.4 0.105 1.4 0.105 0.68 0.135 0.68 0.135 0.56 0.255 0.56 0.255 0.8 0.225 0.8 0.225 1.28 0.485 1.28 0.485 2.13 1.29 2.13 1.29 2.05 2.35 2.05 2.35 1.81 4.275 1.81 4.275 0.8 4.935 0.8 4.935 0.68 5.055 0.68 ;
      POLYGON 2.415 1.45 2.375 1.45 2.375 1.57 2.23 1.57 2.23 1.93 0.905 1.93 0.905 2.01 0.785 2.01 0.785 1.62 0.615 1.62 0.615 0.6 0.735 0.6 0.735 1.5 0.905 1.5 0.905 1.81 2.11 1.81 2.11 1.45 2.255 1.45 2.255 1.33 2.295 1.33 2.295 1.17 2.415 1.17 ;
      POLYGON 1.775 1.69 1.515 1.69 1.515 1.4 1.405 1.4 1.405 1.16 1.515 1.16 1.515 0.6 1.635 0.6 1.635 1.57 1.775 1.57 ;
      POLYGON 1.045 1.38 0.925 1.38 0.925 1.26 0.855 1.26 0.855 0.48 0.495 0.48 0.495 1.16 0.345 1.16 0.345 0.92 0.375 0.92 0.375 0.36 0.975 0.36 0.975 1.14 1.045 1.14 ;
  END
END MX4X4

MACRO MDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX1 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 1.09 0.86 1.425 ;
        RECT 0.65 1.095 0.83 1.435 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.065 0.96 6.185 1.2 ;
        RECT 5.87 0.96 6.185 1.145 ;
        RECT 5.87 0.885 6.02 1.145 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.21 7.625 1.41 ;
        RECT 7.265 1.21 7.525 1.435 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.765 0.97 7.885 1.21 ;
        RECT 7.555 0.94 7.815 1.09 ;
        RECT 6.545 0.97 7.885 1.09 ;
        RECT 6.545 0.97 6.665 1.44 ;
    END
  END S0
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.295 0.265 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.665 -0.18 7.785 0.82 ;
        RECT 6.065 -0.18 6.185 0.64 ;
        RECT 3.795 0.39 4.035 0.51 ;
        RECT 3.795 -0.18 3.915 0.51 ;
        RECT 2.015 -0.18 2.135 0.68 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.445 1.795 7.565 2.79 ;
        RECT 6.065 1.56 6.185 2.79 ;
        RECT 3.795 2.07 4.035 2.19 ;
        RECT 3.795 2.07 3.915 2.79 ;
        RECT 1.715 2.01 1.955 2.13 ;
        RECT 1.715 2.01 1.835 2.79 ;
        RECT 0.565 1.85 0.685 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.205 0.82 8.125 0.82 8.125 1.68 8.045 1.68 8.045 1.8 7.925 1.8 7.925 1.675 6.945 1.675 6.945 1.24 7.065 1.24 7.065 1.555 8.005 1.555 8.005 0.7 8.085 0.7 8.085 0.58 8.205 0.58 ;
      POLYGON 7.145 0.85 6.425 0.85 6.425 1.56 6.825 1.56 6.825 2.21 6.705 2.21 6.705 1.68 6.305 1.68 6.305 1.44 5.355 1.44 5.355 1.59 5.255 1.59 5.255 1.99 5.135 1.99 5.135 1.47 5.235 1.47 5.235 0.72 5.135 0.72 5.135 0.6 5.375 0.6 5.375 0.72 5.355 0.72 5.355 1.32 6.305 1.32 6.305 0.73 7.025 0.73 7.025 0.59 7.145 0.59 ;
      POLYGON 5.765 1.86 5.645 1.86 5.645 1.98 5.495 1.98 5.495 2.23 4.895 2.23 4.895 0.48 4.415 0.48 4.415 0.84 4.535 0.84 4.535 1.1 4.415 1.1 4.415 0.96 4.295 0.96 4.295 0.75 3.555 0.75 3.555 0.48 3.075 0.48 3.075 0.98 3.035 0.98 3.035 1.1 3.015 1.1 3.015 1.27 2.455 1.27 2.455 1.39 2.335 1.39 2.335 1.15 2.895 1.15 2.895 0.86 2.955 0.86 2.955 0.36 3.675 0.36 3.675 0.63 4.295 0.63 4.295 0.36 5.705 0.36 5.705 0.81 5.585 0.81 5.585 0.48 5.015 0.48 5.015 1.11 5.115 1.11 5.115 1.35 5.015 1.35 5.015 2.11 5.375 2.11 5.375 1.86 5.525 1.86 5.525 1.74 5.765 1.74 ;
      POLYGON 4.775 1.99 4.655 1.99 4.655 1.56 3.755 1.56 3.755 1.13 3.875 1.13 3.875 1.44 4.655 1.44 4.655 0.72 4.535 0.72 4.535 0.6 4.775 0.6 ;
      POLYGON 4.595 2.25 4.355 2.25 4.355 1.95 3.255 1.95 3.255 2.23 2.075 2.23 2.075 1.89 1.105 1.89 1.105 2.1 0.985 2.1 0.985 1.29 1.035 1.29 1.035 0.68 1.155 0.68 1.155 1.41 1.105 1.41 1.105 1.77 2.195 1.77 2.195 2.11 3.135 2.11 3.135 1.23 3.275 1.23 3.275 1.11 3.395 1.11 3.395 1.35 3.255 1.35 3.255 1.83 4.475 1.83 4.475 2.13 4.595 2.13 ;
      POLYGON 4.195 1.32 4.055 1.32 4.055 1.01 3.635 1.01 3.635 1.59 3.495 1.59 3.495 1.71 3.375 1.71 3.375 1.47 3.515 1.47 3.515 0.99 3.195 0.99 3.195 0.6 3.435 0.6 3.435 0.87 3.635 0.87 3.635 0.89 4.175 0.89 4.175 1.08 4.195 1.08 ;
      POLYGON 2.835 0.72 2.375 0.72 2.375 1.03 2.215 1.03 2.215 1.51 2.575 1.51 2.575 1.47 2.695 1.47 2.695 1.99 2.575 1.99 2.575 1.63 1.595 1.63 1.595 1.37 1.515 1.37 1.515 1.13 1.715 1.13 1.715 1.51 2.095 1.51 2.095 0.91 2.255 0.91 2.255 0.6 2.835 0.6 ;
      POLYGON 1.975 1.39 1.855 1.39 1.855 1.01 1.395 1.01 1.395 1.53 1.475 1.53 1.475 1.65 1.235 1.65 1.235 1.53 1.275 1.53 1.275 0.56 0.915 0.56 0.915 0.97 0.52 0.97 0.52 1.24 0.4 1.24 0.4 0.85 0.795 0.85 0.795 0.44 1.715 0.44 1.715 0.89 1.975 0.89 ;
  END
END MDFFHQX1

MACRO NOR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X4 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.105 1.26 6.775 1.38 ;
        RECT 6.105 1.23 6.365 1.38 ;
        RECT 6.245 1.14 6.365 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 1.26 5.205 1.38 ;
        RECT 4.915 1.23 5.205 1.38 ;
        RECT 4.915 1.14 5.035 1.38 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.455 1.26 3.355 1.38 ;
        RECT 3.235 1 3.355 1.38 ;
        RECT 2.625 1.23 2.885 1.38 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.435 ;
        RECT 1.535 1 1.655 1.435 ;
        RECT 0.755 1.28 1.67 1.4 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 0.76 6.975 0.88 ;
        RECT 6.855 0.59 6.975 0.88 ;
        RECT 6.825 1.5 6.945 2.01 ;
        RECT 2.13 1.5 6.945 1.62 ;
        RECT 6.015 0.59 6.135 0.88 ;
        RECT 5.985 1.5 6.105 2.01 ;
        RECT 5.175 0.59 5.295 0.88 ;
        RECT 4.335 0.59 4.455 0.88 ;
        RECT 3.495 0.59 3.615 0.88 ;
        RECT 2.655 0.59 2.775 0.88 ;
        RECT 2.13 0.76 2.25 1.62 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.815 0.59 1.935 0.88 ;
        RECT 0.975 0.59 1.095 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 7.275 -0.18 7.395 0.64 ;
        RECT 6.435 -0.18 6.555 0.64 ;
        RECT 5.595 -0.18 5.715 0.64 ;
        RECT 4.755 -0.18 4.875 0.64 ;
        RECT 3.915 -0.18 4.035 0.64 ;
        RECT 3.075 -0.18 3.195 0.64 ;
        RECT 2.235 -0.18 2.355 0.64 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 1.335 1.98 1.575 2.15 ;
        RECT 1.335 1.98 1.455 2.79 ;
        RECT 0.495 1.98 0.735 2.15 ;
        RECT 0.495 1.98 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.365 2.25 5.565 2.25 5.565 1.86 4.845 1.86 4.845 2.01 4.725 2.01 4.725 1.86 4.005 1.86 4.005 2.01 3.885 2.01 3.885 1.74 5.685 1.74 5.685 2.13 6.405 2.13 6.405 1.74 6.525 1.74 6.525 2.13 7.245 2.13 7.245 1.56 7.365 1.56 ;
      POLYGON 5.325 2.15 5.205 2.15 5.205 2.25 2.295 2.25 2.295 2.15 2.175 2.15 2.175 1.98 2.415 1.98 2.415 2.13 3.015 2.13 3.015 1.98 3.255 1.98 3.255 2.13 4.245 2.13 4.245 1.98 4.485 1.98 4.485 2.13 5.085 2.13 5.085 1.98 5.325 1.98 ;
      POLYGON 3.615 2.01 3.495 2.01 3.495 1.86 2.775 1.86 2.775 2.01 2.655 2.01 2.655 1.86 1.935 1.86 1.935 2.21 1.815 2.21 1.815 1.86 1.095 1.86 1.095 2.21 0.975 2.21 0.975 1.86 0.255 1.86 0.255 2.21 0.135 2.21 0.135 1.56 0.255 1.56 0.255 1.74 0.975 1.74 0.975 1.56 1.095 1.56 1.095 1.74 1.815 1.74 1.815 1.56 1.935 1.56 1.935 1.74 3.615 1.74 ;
  END
END NOR4X4

MACRO DFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX4 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 0.59 1.515 1.99 ;
        RECT 0.555 1.025 1.515 1.145 ;
        RECT 0.555 0.885 0.8 1.145 ;
        RECT 0.555 0.59 0.675 1.99 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.905 0.94 3.175 1.2 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.18 10.715 1.45 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.615 0.94 11.875 1.155 ;
        RECT 11.615 0.94 11.735 1.32 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.235 2.13 8.475 2.25 ;
        RECT 7.595 2.01 8.355 2.13 ;
        RECT 7.595 1.7 7.715 2.13 ;
        RECT 6.995 1.7 7.715 1.82 ;
        RECT 5.795 2.13 7.115 2.25 ;
        RECT 6.995 1.7 7.115 2.25 ;
        RECT 5.795 1.52 5.915 2.25 ;
        RECT 5.235 1.52 5.915 1.64 ;
        RECT 5.235 1.52 5.495 1.67 ;
        RECT 5.065 1.43 5.355 1.55 ;
    END
  END SN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.865 -0.18 11.985 0.82 ;
        RECT 10.515 -0.18 10.635 0.78 ;
        RECT 9.115 -0.18 9.235 0.64 ;
        RECT 5.205 -0.18 5.445 0.34 ;
        RECT 2.595 0.46 2.835 0.58 ;
        RECT 2.715 -0.18 2.835 0.58 ;
        RECT 1.815 -0.18 1.935 0.64 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.865 1.46 11.985 2.79 ;
        RECT 10.675 1.84 10.795 2.79 ;
        RECT 8.595 2.01 8.835 2.13 ;
        RECT 8.595 2.01 8.715 2.79 ;
        RECT 7.355 1.94 7.475 2.79 ;
        RECT 7.235 1.94 7.475 2.06 ;
        RECT 5.045 2.27 5.285 2.79 ;
        RECT 3.785 2.04 3.905 2.79 ;
        RECT 3.665 2.04 3.905 2.16 ;
        RECT 2.655 1.56 2.775 2.79 ;
        RECT 1.815 1.44 1.935 2.79 ;
        RECT 0.975 1.34 1.095 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.625 1.56 11.375 1.56 11.375 0.7 11.445 0.7 11.445 0.48 10.875 0.48 10.875 0.94 11.015 0.94 11.015 1.06 10.755 1.06 10.755 1.04 10.195 1.04 10.195 1.16 10.075 1.16 10.075 2.25 9.475 2.25 9.475 1.89 7.835 1.89 7.835 1.58 6.875 1.58 6.875 2.01 6.275 2.01 6.275 0.98 6.395 0.98 6.395 0.49 5.915 0.49 5.915 1.07 5.675 1.07 5.675 0.95 5.795 0.95 5.795 0.37 6.515 0.37 6.515 1.1 6.395 1.1 6.395 1.89 6.755 1.89 6.755 1.46 7.955 1.46 7.955 1.77 9.425 1.77 9.425 1.54 9.355 1.54 9.355 1.42 9.595 1.42 9.595 1.54 9.545 1.54 9.545 1.77 9.595 1.77 9.595 2.13 9.955 2.13 9.955 0.92 10.755 0.92 10.755 0.36 11.565 0.36 11.565 0.82 11.495 0.82 11.495 1.44 11.625 1.44 ;
      POLYGON 11.255 1.69 11.215 1.69 11.215 2.08 11.095 2.08 11.095 1.69 10.195 1.69 10.195 1.34 10.315 1.34 10.315 1.57 11.135 1.57 11.135 0.72 10.995 0.72 10.995 0.6 11.255 0.6 ;
      POLYGON 9.995 0.74 9.835 0.74 9.835 2.01 9.715 2.01 9.715 0.74 9.475 0.74 9.475 0.88 8.795 0.88 8.795 1 8.555 1 8.555 0.88 8.675 0.88 8.675 0.76 9.355 0.76 9.355 0.62 9.875 0.62 9.875 0.5 9.995 0.5 ;
      POLYGON 9.595 1.24 8.315 1.24 8.315 1.1 6.875 1.1 6.875 0.98 8.435 0.98 8.435 1.12 9.355 1.12 9.355 1.1 9.595 1.1 ;
      POLYGON 9.235 1.54 8.335 1.54 8.335 1.65 8.075 1.65 8.075 1.34 6.635 1.34 6.635 1.77 6.515 1.77 6.515 1.22 6.635 1.22 6.635 0.55 6.755 0.55 6.755 0.74 7.875 0.74 7.875 0.6 8.115 0.6 8.115 0.72 7.995 0.72 7.995 0.86 6.755 0.86 6.755 1.22 8.195 1.22 8.195 1.42 9.235 1.42 ;
      POLYGON 8.475 0.68 8.355 0.68 8.355 0.48 7.755 0.48 7.755 0.62 7.455 0.62 7.455 0.5 7.635 0.5 7.635 0.36 8.475 0.36 ;
      POLYGON 6.275 0.73 6.155 0.73 6.155 1.97 6.035 1.97 6.035 1.31 4.945 1.31 4.945 1.57 4.445 1.57 4.445 1.92 2.895 1.92 2.895 1.44 2.515 1.44 2.515 1.12 2.635 1.12 2.635 1.32 3.015 1.32 3.015 1.8 4.325 1.8 4.325 1.45 4.825 1.45 4.825 1.19 6.035 1.19 6.035 0.61 6.275 0.61 ;
      POLYGON 5.675 0.73 5.435 0.73 5.435 0.58 4.965 0.58 4.965 0.48 4.425 0.48 4.425 0.62 4.185 0.62 4.185 0.5 4.305 0.5 4.305 0.36 5.085 0.36 5.085 0.46 5.555 0.46 5.555 0.61 5.675 0.61 ;
      POLYGON 5.675 1.91 4.685 1.91 4.685 1.97 4.565 1.97 4.565 1.69 4.685 1.69 4.685 1.79 5.675 1.79 ;
      POLYGON 5.675 2.25 5.405 2.25 5.405 2.15 4.925 2.15 4.925 2.21 4.795 2.21 4.795 2.25 4.025 2.25 4.025 2.13 4.675 2.13 4.675 2.09 4.805 2.09 4.805 2.03 5.525 2.03 5.525 2.13 5.675 2.13 ;
      POLYGON 4.845 0.72 4.705 0.72 4.705 1.28 3.705 1.28 3.705 0.72 3.585 0.72 3.585 0.6 3.825 0.6 3.825 1.16 4.585 1.16 4.585 0.6 4.845 0.6 ;
      POLYGON 4.465 1.04 4.225 1.04 4.225 0.86 3.945 0.86 3.945 0.48 3.075 0.48 3.075 0.82 2.355 0.82 2.355 1.56 2.415 1.56 2.415 1.9 2.175 1.9 2.175 1.56 2.235 1.56 2.235 1.2 1.635 1.2 1.635 1.08 2.235 1.08 2.235 0.5 2.355 0.5 2.355 0.7 2.955 0.7 2.955 0.36 4.065 0.36 4.065 0.74 4.345 0.74 4.345 0.92 4.465 0.92 ;
      POLYGON 3.585 1.3 3.415 1.3 3.415 1.44 3.255 1.44 3.255 1.68 3.135 1.68 3.135 1.32 3.295 1.32 3.295 0.72 3.195 0.72 3.195 0.6 3.435 0.6 3.435 0.72 3.415 0.72 3.415 1.18 3.585 1.18 ;
  END
END DFFSRHQX4

MACRO NAND4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX2 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.035 1.21 4.335 1.44 ;
        RECT 4.075 1.185 4.335 1.44 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.26 3.315 1.435 ;
        RECT 2.915 1.23 3.175 1.435 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.18 2.595 1.45 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 1.22 0.565 1.38 ;
        RECT 0.175 1.12 0.415 1.25 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9696 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.195 0.65 4.435 0.77 ;
        RECT 2.095 0.94 4.315 1.06 ;
        RECT 4.195 0.65 4.315 1.06 ;
        RECT 3.935 1.56 4.055 2.21 ;
        RECT 1.415 1.57 4.055 1.69 ;
        RECT 3.095 1.56 3.215 2.21 ;
        RECT 2.255 1.57 2.375 2.21 ;
        RECT 2.1 1.57 2.375 2.015 ;
        RECT 2.095 0.94 2.215 1.69 ;
        RECT 1.415 1.56 1.535 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 1.345 -0.18 1.465 0.64 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 4.355 1.56 4.475 2.79 ;
        RECT 3.515 1.81 3.635 2.79 ;
        RECT 2.675 1.81 2.795 2.79 ;
        RECT 1.835 1.81 1.955 2.79 ;
        RECT 0.995 1.77 1.115 2.79 ;
        RECT 0.265 1.5 0.385 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.795 0.65 4.675 0.65 4.675 0.53 3.955 0.53 3.955 0.65 3.835 0.65 3.835 0.53 3.175 0.53 3.175 0.58 2.935 0.58 2.935 0.46 3.055 0.46 3.055 0.41 4.795 0.41 ;
      POLYGON 3.595 0.77 3.475 0.77 3.475 0.82 2.245 0.82 2.245 0.77 2.125 0.77 2.125 0.65 2.365 0.65 2.365 0.7 3.355 0.7 3.355 0.65 3.595 0.65 ;
      POLYGON 2.785 0.58 2.545 0.58 2.545 0.53 1.885 0.53 1.885 0.88 0.925 0.88 0.925 0.59 1.045 0.59 1.045 0.76 1.765 0.76 1.765 0.41 2.665 0.41 2.665 0.46 2.785 0.46 ;
      POLYGON 1.335 1.32 0.805 1.32 0.805 1.62 0.685 1.62 0.685 1.1 0.535 1.1 0.535 0.68 0.655 0.68 0.655 0.98 0.805 0.98 0.805 1.2 1.335 1.2 ;
  END
END NAND4BX2

MACRO AO22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.935 0.99 1.055 1.23 ;
        RECT 0.65 0.99 1.055 1.11 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.315 0.89 1.435 1.255 ;
        RECT 1.175 0.89 1.435 1.1 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.985 0.415 1.44 ;
        RECT 0.295 0.965 0.415 1.44 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 1.02 1.96 1.44 ;
        RECT 1.795 1 1.915 1.44 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.665 1.145 2.785 2.21 ;
        RECT 2.42 1.145 2.785 1.265 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.375 0.59 2.495 1.025 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.795 -0.18 2.915 0.64 ;
        RECT 1.955 -0.18 2.075 0.64 ;
        RECT 0.41 -0.18 0.53 0.83 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 3.085 1.56 3.205 2.79 ;
        RECT 2.185 2.01 2.425 2.15 ;
        RECT 2.185 2.01 2.305 2.79 ;
        RECT 0.615 2.08 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.255 1.15 2.135 1.15 2.135 0.88 1.675 0.88 1.675 1.56 1.695 1.56 1.695 1.68 1.455 1.68 1.455 1.56 1.555 1.56 1.555 0.77 1.035 0.77 1.035 0.65 1.675 0.65 1.675 0.76 2.255 0.76 ;
      POLYGON 2.055 1.92 1.095 1.92 1.095 1.68 0.075 1.68 0.075 1.56 1.215 1.56 1.215 1.8 1.935 1.8 1.935 1.56 2.055 1.56 ;
  END
END AO22X2

MACRO BUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.87 0.825 3.99 1.305 ;
        RECT 3.84 0.825 3.99 1.28 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.69 0.715 2.93 0.835 ;
        RECT 2.75 1.295 2.87 2.21 ;
        RECT 0.23 0.76 2.81 0.88 ;
        RECT 2.57 1.295 2.87 1.415 ;
        RECT 0.23 1.27 2.69 1.39 ;
        RECT 1.85 0.71 2.09 0.88 ;
        RECT 1.91 1.27 2.03 2.21 ;
        RECT 1.01 0.71 1.25 0.88 ;
        RECT 1.07 1.27 1.19 2.21 ;
        RECT 0.36 0.76 0.51 1.145 ;
        RECT 0.36 0.76 0.48 1.39 ;
        RECT 0.23 1.27 0.35 2.21 ;
        RECT 0.23 0.64 0.35 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 4.01 -0.18 4.13 0.705 ;
        RECT 3.17 -0.18 3.29 0.705 ;
        RECT 2.33 -0.18 2.45 0.64 ;
        RECT 1.49 -0.18 1.61 0.64 ;
        RECT 0.65 -0.18 0.77 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 4.01 1.465 4.13 2.79 ;
        RECT 3.17 1.465 3.29 2.79 ;
        RECT 2.33 1.51 2.45 2.79 ;
        RECT 1.49 1.51 1.61 2.79 ;
        RECT 0.65 1.51 0.77 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.71 2.115 3.59 2.115 3.59 1.15 3.19 1.15 3.19 1.175 2.95 1.175 2.95 1.15 0.87 1.15 0.87 1.03 3.59 1.03 3.59 0.655 3.71 0.655 ;
  END
END BUFX8

MACRO DFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX1 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.455 0.915 1.725 ;
        RECT 0.65 1.44 0.8 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.985 1.49 5.225 1.725 ;
        RECT 4.945 1.495 5.205 1.75 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 2.205 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.185 0.68 5.425 0.8 ;
        RECT 5.185 -0.18 5.305 0.8 ;
        RECT 3.625 0.45 3.865 0.57 ;
        RECT 3.745 -0.18 3.865 0.57 ;
        RECT 1.925 -0.18 2.045 0.86 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.185 1.87 5.305 2.79 ;
        RECT 3.525 2.29 3.765 2.79 ;
        RECT 1.805 2.29 2.045 2.79 ;
        RECT 0.555 1.845 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.805 1.61 5.725 1.61 5.725 1.99 5.605 1.99 5.605 1.49 5.685 1.49 5.685 1.04 4.87 1.04 4.87 0.5 4.105 0.5 4.105 0.81 3.385 0.81 3.385 0.5 3.025 0.5 3.025 1.17 3.225 1.17 3.225 1.29 2.665 1.29 2.665 1.53 2.585 1.53 2.585 1.65 2.465 1.65 2.465 1.41 2.545 1.41 2.545 1.17 2.905 1.17 2.905 0.38 3.505 0.38 3.505 0.69 3.985 0.69 3.985 0.38 4.265 0.38 4.265 0.36 4.505 0.36 4.505 0.38 4.99 0.38 4.99 0.92 5.665 0.92 5.665 0.62 5.785 0.62 5.785 0.74 5.805 0.74 ;
      POLYGON 5.565 1.37 4.805 1.37 4.805 1.41 4.705 1.41 4.705 2.17 2.925 2.17 2.925 2.25 2.275 2.25 2.275 2.17 0.975 2.17 0.975 1.845 1.035 1.845 1.035 0.68 1.155 0.68 1.155 2.05 2.395 2.05 2.395 2.13 2.805 2.13 2.805 1.61 2.785 1.61 2.785 1.49 3.025 1.49 3.025 1.61 2.925 1.61 2.925 2.05 4.585 2.05 4.585 1.65 4.125 1.65 4.125 1.41 4.245 1.41 4.245 1.53 4.585 1.53 4.585 1.25 4.685 1.25 4.685 1.17 4.805 1.17 4.805 1.25 5.565 1.25 ;
      POLYGON 4.725 1.05 4.005 1.05 4.005 1.77 4.345 1.77 4.345 1.81 4.465 1.81 4.465 1.93 4.225 1.93 4.225 1.89 3.885 1.89 3.885 1.45 3.705 1.45 3.705 1.57 3.585 1.57 3.585 1.33 3.885 1.33 3.885 0.93 4.605 0.93 4.605 0.62 4.725 0.62 ;
      POLYGON 3.765 1.21 3.465 1.21 3.465 1.93 3.045 1.93 3.045 1.81 3.345 1.81 3.345 1.05 3.145 1.05 3.145 0.62 3.265 0.62 3.265 0.93 3.465 0.93 3.465 1.09 3.645 1.09 3.645 0.97 3.765 0.97 ;
      POLYGON 2.785 0.8 2.345 0.8 2.345 1.77 2.685 1.77 2.685 2.01 2.565 2.01 2.565 1.89 2.225 1.89 2.225 1.53 1.645 1.53 1.645 1.41 2.225 1.41 2.225 0.68 2.785 0.68 ;
      POLYGON 2.105 1.2 1.525 1.2 1.525 1.81 1.565 1.81 1.565 1.93 1.325 1.93 1.325 1.81 1.405 1.81 1.405 0.74 1.425 0.74 1.425 0.56 0.915 0.56 0.915 0.97 0.535 0.97 0.535 1.24 0.415 1.24 0.415 0.85 0.795 0.85 0.795 0.44 1.545 0.44 1.545 0.86 1.525 0.86 1.525 1.08 2.105 1.08 ;
  END
END DFFQX1

MACRO DFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX1 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.725 1.19 2.015 1.38 ;
        RECT 1.655 1.17 1.925 1.33 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.97 2.13 6.475 2.25 ;
        RECT 5.97 1.76 6.09 2.25 ;
        RECT 5.215 1.76 6.09 1.88 ;
        RECT 3.745 2.13 5.335 2.25 ;
        RECT 5.215 1.76 5.335 2.25 ;
        RECT 3.745 1.7 3.865 2.25 ;
        RECT 3.1 1.7 3.865 1.82 ;
        RECT 2.305 1.89 3.22 2.01 ;
        RECT 3.1 1.7 3.22 2.01 ;
        RECT 2.305 1.175 2.54 1.435 ;
        RECT 2.255 1.17 2.495 1.29 ;
        RECT 2.305 1.17 2.425 2.01 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.575 1.23 8.975 1.38 ;
        RECT 8.575 1.21 8.715 1.45 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.875 1.175 10.135 1.38 ;
        RECT 9.875 1.03 9.995 1.38 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 10.115 -0.18 10.235 0.91 ;
        RECT 8.735 -0.18 8.855 0.85 ;
        RECT 7.155 -0.18 7.275 0.68 ;
        RECT 1.975 -0.18 2.095 0.81 ;
        RECT 0.555 -0.18 0.675 0.82 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 10.115 1.5 10.235 2.79 ;
        RECT 8.675 1.81 8.795 2.79 ;
        RECT 7.215 1.93 7.335 2.79 ;
        RECT 7.095 1.93 7.335 2.05 ;
        RECT 5.575 2 5.695 2.79 ;
        RECT 5.455 2 5.695 2.12 ;
        RECT 3.385 1.94 3.625 2.06 ;
        RECT 3.385 1.94 3.505 2.79 ;
        RECT 1.825 1.74 1.945 2.79 ;
        RECT 1.705 1.74 1.945 1.86 ;
        RECT 0.555 1.69 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.875 1.62 9.635 1.62 9.635 0.79 9.695 0.79 9.695 0.56 9.095 0.56 9.095 1.09 8.455 1.09 8.455 1.13 8.195 1.13 8.195 1.01 8.335 1.01 8.335 0.48 7.715 0.48 7.715 1.21 7.835 1.21 7.835 1.33 7.595 1.33 7.595 0.92 6.295 0.92 6.295 1.16 5.035 1.16 5.035 1.04 6.175 1.04 6.175 0.8 7.595 0.8 7.595 0.36 8.455 0.36 8.455 0.97 8.975 0.97 8.975 0.44 9.015 0.44 9.015 0.36 9.255 0.36 9.255 0.44 9.815 0.44 9.815 0.91 9.755 0.91 9.755 1.5 9.875 1.5 ;
      POLYGON 9.455 1.33 9.215 1.33 9.215 2.05 9.095 2.05 9.095 1.69 8.315 1.69 8.315 2.25 7.455 2.25 7.455 1.81 6.975 1.81 6.975 2.01 6.255 2.01 6.255 1.64 5.095 1.64 5.095 2.01 4.015 2.01 4.015 1.06 4.135 1.06 4.135 1.89 4.495 1.89 4.495 1.04 4.555 1.04 4.555 0.84 4.675 0.84 4.675 1.16 4.615 1.16 4.615 1.89 4.975 1.89 4.975 1.52 6.375 1.52 6.375 1.89 6.855 1.89 6.855 1.69 7.575 1.69 7.575 2.13 8.195 2.13 8.195 1.31 8.315 1.31 8.315 1.57 9.095 1.57 9.095 1.21 9.215 1.21 9.215 0.68 9.455 0.68 ;
      POLYGON 8.215 0.72 8.075 0.72 8.075 1.69 8.055 1.69 8.055 2.01 7.935 2.01 7.935 1.57 7.355 1.57 7.355 1.16 6.415 1.16 6.415 1.04 7.475 1.04 7.475 1.45 7.955 1.45 7.955 0.6 8.215 0.6 ;
      POLYGON 7.235 1.4 6.735 1.4 6.735 1.77 6.495 1.77 6.495 1.65 6.615 1.65 6.615 1.4 4.855 1.4 4.855 1.77 4.735 1.77 4.735 1.28 4.795 1.28 4.795 0.5 4.915 0.5 4.915 0.74 5.815 0.74 5.815 0.6 6.055 0.6 6.055 0.72 5.935 0.72 5.935 0.86 4.915 0.86 4.915 1.28 7.235 1.28 ;
      POLYGON 6.415 0.68 6.295 0.68 6.295 0.48 5.635 0.48 5.635 0.62 5.395 0.62 5.395 0.5 5.515 0.5 5.515 0.36 6.415 0.36 ;
      POLYGON 4.435 0.92 4.375 0.92 4.375 1.77 4.255 1.77 4.255 0.94 3.895 0.94 3.895 1.23 2.66 1.23 2.66 1.05 1.735 1.05 1.735 0.51 0.915 0.51 0.915 1.24 0.795 1.24 0.795 0.39 1.855 0.39 1.855 0.93 2.78 0.93 2.78 1.11 3.775 1.11 3.775 0.82 4.255 0.82 4.255 0.8 4.315 0.8 4.315 0.5 4.435 0.5 ;
      POLYGON 4.075 0.68 3.955 0.68 3.955 0.7 3.655 0.7 3.655 0.99 2.9 0.99 2.9 0.81 2.755 0.81 2.755 0.69 3.02 0.69 3.02 0.87 3.535 0.87 3.535 0.58 3.835 0.58 3.835 0.56 4.075 0.56 ;
      POLYGON 3.895 1.58 2.785 1.58 2.785 1.77 2.545 1.77 2.545 1.555 2.665 1.555 2.665 1.46 3.895 1.46 ;
      POLYGON 3.415 0.75 3.175 0.75 3.175 0.57 2.515 0.57 2.515 0.81 2.395 0.81 2.395 0.45 3.295 0.45 3.295 0.63 3.415 0.63 ;
      POLYGON 3.265 2.25 2.065 2.25 2.065 1.62 1.405 1.62 1.405 1.67 1.285 1.67 1.285 0.63 1.615 0.63 1.615 0.75 1.405 0.75 1.405 1.5 2.185 1.5 2.185 2.13 3.265 2.13 ;
      POLYGON 1.705 2.25 0.975 2.25 0.975 1.82 1.035 1.82 1.035 1.48 0.415 1.48 0.415 1.24 0.535 1.24 0.535 1.36 1.035 1.36 1.035 0.68 1.155 0.68 1.155 1.94 1.095 1.94 1.095 2.13 1.705 2.13 ;
  END
END DFFSRHQX1

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.855 1.28 0.975 1.56 ;
        RECT 0.68 1.44 0.975 1.56 ;
        RECT 0.65 1.465 0.8 1.725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 1.18 2.835 1.3 ;
        RECT 2.045 1.18 2.305 1.38 ;
        RECT 1.915 1.14 2.155 1.3 ;
        RECT 1.335 1.36 1.575 1.48 ;
        RECT 1.455 1.18 1.575 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.295 0.29 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.395 -0.18 2.515 0.78 ;
        RECT 0.495 0.55 0.735 0.67 ;
        RECT 0.615 -0.18 0.735 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.275 1.74 2.395 2.79 ;
        RECT 0.59 2.16 0.83 2.28 ;
        RECT 0.59 2.16 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.075 1.74 2.815 1.74 2.815 1.86 2.695 1.86 2.695 1.62 1.955 1.62 1.955 2.24 1.715 2.24 1.715 2.12 1.835 2.12 1.835 1.5 2.815 1.5 2.815 1.62 2.955 1.62 2.955 0.78 2.815 0.78 2.815 0.54 2.935 0.54 2.935 0.66 3.075 0.66 ;
      POLYGON 2.515 1.06 2.275 1.06 2.275 1.02 1.215 1.02 1.215 1.68 1.31 1.68 1.31 1.8 1.07 1.8 1.07 1.68 1.095 1.68 1.095 0.6 1.335 0.6 1.335 0.72 1.215 0.72 1.215 0.9 2.395 0.9 2.395 0.94 2.515 0.94 ;
      POLYGON 1.875 0.78 1.755 0.78 1.755 0.48 0.975 0.48 0.975 1.16 0.55 1.16 0.55 1.28 0.53 1.28 0.53 1.92 1.475 1.92 1.475 1.86 1.55 1.86 1.55 1.74 1.67 1.74 1.67 1.98 1.595 1.98 1.595 2.04 0.41 2.04 0.41 1.04 0.855 1.04 0.855 0.36 1.875 0.36 ;
  END
END XOR2X1

MACRO NAND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X4 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.585 1.08 6.825 1.2 ;
        RECT 5.865 1.26 6.705 1.38 ;
        RECT 6.585 1.08 6.705 1.38 ;
        RECT 6.105 1.23 6.365 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.505 1.08 5.745 1.2 ;
        RECT 4.135 1.26 5.625 1.38 ;
        RECT 5.505 1.08 5.625 1.38 ;
        RECT 5.235 1.23 5.625 1.38 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.455 1.26 3.035 1.38 ;
        RECT 2.625 1.23 2.885 1.38 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.26 1.315 1.38 ;
        RECT 0.885 1.23 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9392 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.265 0.84 7.025 0.96 ;
        RECT 6.905 0.64 7.025 0.96 ;
        RECT 6.435 1.5 6.555 2.21 ;
        RECT 0.555 1.5 6.555 1.62 ;
        RECT 6.065 0.64 6.185 0.96 ;
        RECT 5.595 1.5 5.715 2.21 ;
        RECT 2.215 0.99 5.385 1.11 ;
        RECT 5.265 0.84 5.385 1.11 ;
        RECT 4.755 1.5 4.875 2.21 ;
        RECT 3.915 1.5 4.035 2.21 ;
        RECT 3.075 1.5 3.195 2.21 ;
        RECT 2.235 1.5 2.355 2.21 ;
        RECT 2.1 1.465 2.335 1.725 ;
        RECT 2.215 0.99 2.335 1.725 ;
        RECT 1.395 1.5 1.515 2.21 ;
        RECT 0.555 1.5 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 1.395 -0.18 1.515 0.69 ;
        RECT 0.555 -0.18 0.675 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.855 1.56 6.975 2.79 ;
        RECT 6.015 1.74 6.135 2.79 ;
        RECT 5.175 1.74 5.295 2.79 ;
        RECT 4.335 1.74 4.455 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.445 0.69 7.325 0.69 7.325 0.48 6.605 0.48 6.605 0.69 6.485 0.69 6.485 0.48 5.765 0.48 5.765 0.69 5.645 0.69 5.645 0.48 4.905 0.48 4.905 0.63 4.665 0.63 4.665 0.48 4.065 0.48 4.065 0.63 3.825 0.63 3.825 0.51 3.945 0.51 3.945 0.36 7.445 0.36 ;
      POLYGON 5.405 0.72 5.145 0.72 5.145 0.87 2.355 0.87 2.355 0.82 2.175 0.82 2.175 0.7 2.475 0.7 2.475 0.75 3.075 0.75 3.075 0.63 3.195 0.63 3.195 0.75 4.305 0.75 4.305 0.63 4.425 0.63 4.425 0.75 5.025 0.75 5.025 0.6 5.405 0.6 ;
      POLYGON 3.675 0.63 3.435 0.63 3.435 0.51 2.835 0.51 2.835 0.63 2.595 0.63 2.595 0.51 1.935 0.51 1.935 0.93 0.135 0.93 0.135 0.64 0.255 0.64 0.255 0.81 0.975 0.81 0.975 0.64 1.095 0.64 1.095 0.81 1.815 0.81 1.815 0.39 3.555 0.39 3.555 0.51 3.675 0.51 ;
  END
END NAND4X4

MACRO AOI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.095 1.96 1.435 ;
        RECT 1.78 0.98 1.9 1.32 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.41 1.38 1.725 ;
        RECT 1.24 1.22 1.36 1.725 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.34 0.98 1.46 ;
        RECT 0.86 1.22 0.98 1.46 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.34 0.8 1.725 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3196 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.69 0.84 0.81 ;
        RECT 0.24 0.74 0.72 0.86 ;
        RECT 0.38 1.27 0.5 2.21 ;
        RECT 0.24 1.27 0.5 1.39 ;
        RECT 0.24 0.74 0.36 1.39 ;
        RECT 0.07 0.885 0.36 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.92 -0.18 2.04 0.86 ;
        RECT 1.08 -0.18 1.2 0.86 ;
        RECT 0.18 0.5 0.42 0.62 ;
        RECT 0.18 -0.18 0.3 0.62 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.02 1.845 1.14 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.9 1.74 1.5 1.74 1.5 1.1 0.74 1.1 0.74 1.15 0.48 1.15 0.48 1.03 0.62 1.03 0.62 0.98 1.5 0.98 1.5 0.62 1.62 0.62 1.62 1.62 1.9 1.62 ;
  END
END AOI2BB1X1

MACRO AOI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X4 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 1.04 3.32 1.16 ;
        RECT 0.65 1.04 0.8 1.435 ;
    END
  END B0
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.13 0.985 4.28 1.44 ;
        RECT 4.13 0.965 4.25 1.44 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 0.78 3.7 1.235 ;
        RECT 3.58 0.76 3.7 1.235 ;
    END
  END A0N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9664 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.18 0.76 3.2 0.88 ;
        RECT 3.08 0.59 3.2 0.88 ;
        RECT 2.26 1.595 2.38 2.21 ;
        RECT 2.24 0.59 2.36 0.88 ;
        RECT 0.18 1.595 2.38 1.715 ;
        RECT 1.4 0.59 1.52 0.88 ;
        RECT 0.98 1.56 1.1 2.21 ;
        RECT 0.56 0.59 0.68 0.88 ;
        RECT 0.305 1.595 0.565 1.96 ;
        RECT 0.18 1.595 0.565 1.93 ;
        RECT 0.18 0.76 0.3 1.93 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 4.34 -0.18 4.46 0.64 ;
        RECT 3.5 -0.18 3.62 0.64 ;
        RECT 2.66 -0.18 2.78 0.64 ;
        RECT 1.82 -0.18 1.94 0.64 ;
        RECT 0.98 -0.18 1.1 0.64 ;
        RECT 0.14 -0.18 0.26 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.3 1.595 3.42 2.79 ;
        RECT 1.62 1.835 1.74 2.79 ;
        RECT 0.22 2.08 0.46 2.2 ;
        RECT 0.22 2.08 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.06 2.21 3.94 2.21 3.94 1.68 3.89 1.68 3.89 1.475 1.22 1.475 1.22 1.4 1.08 1.4 1.08 1.28 1.34 1.28 1.34 1.355 2.32 1.355 2.32 1.3 2.56 1.3 2.56 1.355 3.89 1.355 3.89 0.725 3.92 0.725 3.92 0.59 4.04 0.59 4.04 0.845 4.01 0.845 4.01 1.56 4.06 1.56 ;
  END
END AOI2BB1X4

MACRO CLKINVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX16 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.728 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.205 5.495 1.325 ;
        RECT 0.885 1.205 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.5 5.735 1.62 ;
        RECT 5.615 0.79 5.735 1.62 ;
        RECT 5.58 1.465 5.73 1.725 ;
        RECT 5.595 1.465 5.715 2.21 ;
        RECT 0.615 0.79 5.735 0.91 ;
        RECT 5.595 0.67 5.715 0.91 ;
        RECT 4.695 0.74 4.935 0.91 ;
        RECT 4.755 1.47 4.875 2.21 ;
        RECT 3.855 0.74 4.095 0.91 ;
        RECT 3.915 1.47 4.035 2.21 ;
        RECT 3.015 0.74 3.255 0.91 ;
        RECT 3.075 1.465 3.195 2.21 ;
        RECT 2.175 0.74 2.415 0.91 ;
        RECT 2.235 1.465 2.355 2.21 ;
        RECT 1.335 0.74 1.575 0.91 ;
        RECT 1.395 1.465 1.515 2.21 ;
        RECT 0.495 0.74 0.735 0.86 ;
        RECT 0.555 1.465 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 6.015 -0.18 6.135 0.67 ;
        RECT 5.175 -0.18 5.295 0.67 ;
        RECT 4.335 -0.18 4.455 0.67 ;
        RECT 3.495 -0.18 3.615 0.67 ;
        RECT 2.655 -0.18 2.775 0.67 ;
        RECT 1.815 -0.18 1.935 0.67 ;
        RECT 0.975 -0.18 1.095 0.665 ;
        RECT 0.135 -0.18 0.255 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 6.015 1.47 6.135 2.79 ;
        RECT 5.175 1.74 5.295 2.79 ;
        RECT 4.335 1.74 4.455 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
END CLKINVX16

MACRO MXI2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X8 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.555 1.27 1.675 ;
        RECT 1.15 1.405 1.27 1.675 ;
        RECT 0.41 1.505 0.53 1.745 ;
        RECT 0.36 1.465 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.95 1.415 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.95 1.175 2.25 1.405 ;
        RECT 1.95 1.165 2.07 1.405 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.79 1.22 5.91 2.2 ;
        RECT 4.17 0.79 5.91 0.91 ;
        RECT 5.79 0.67 5.91 0.91 ;
        RECT 3.26 1.22 5.91 1.34 ;
        RECT 5.48 0.79 5.6 1.34 ;
        RECT 4.89 0.74 5.13 0.91 ;
        RECT 4.95 1.22 5.07 2.2 ;
        RECT 4.05 0.74 4.29 0.86 ;
        RECT 4.11 1.22 4.23 2.205 ;
        RECT 3.26 1.175 3.41 1.435 ;
        RECT 3.27 0.68 3.39 2.205 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.37 -0.18 5.49 0.67 ;
        RECT 4.53 -0.18 4.65 0.67 ;
        RECT 3.69 -0.18 3.81 0.67 ;
        RECT 2.85 -0.18 2.97 0.73 ;
        RECT 2.01 -0.18 2.13 0.805 ;
        RECT 0.67 -0.18 0.79 0.805 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.37 1.46 5.49 2.79 ;
        RECT 4.53 1.46 4.65 2.79 ;
        RECT 3.69 1.46 3.81 2.79 ;
        RECT 2.85 1.555 2.97 2.79 ;
        RECT 2.01 1.555 2.13 2.79 ;
        RECT 0.67 1.965 0.79 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.14 1.32 2.73 1.32 2.73 1.675 2.55 1.675 2.55 2.205 2.43 2.205 2.43 1.555 2.61 1.555 2.61 0.805 2.43 0.805 2.43 0.565 2.55 0.565 2.55 0.685 2.73 0.685 2.73 1.2 3.14 1.2 ;
      POLYGON 2.49 1.24 2.37 1.24 2.37 1.045 1.83 1.045 1.83 1.985 1.49 1.985 1.49 2.025 1.25 2.025 1.25 1.905 1.37 1.905 1.37 1.865 1.71 1.865 1.71 1.045 1.39 1.045 1.39 0.805 1.31 0.805 1.31 0.565 1.43 0.565 1.43 0.685 1.51 0.685 1.51 0.925 2.49 0.925 ;
      POLYGON 1.59 1.745 1.47 1.745 1.47 1.285 1.15 1.285 1.15 1.055 0.24 1.055 0.24 1.845 0.29 1.845 0.29 2.085 0.17 2.085 0.17 1.965 0.12 1.965 0.12 0.685 0.25 0.685 0.25 0.565 0.37 0.565 0.37 0.805 0.24 0.805 0.24 0.935 1.15 0.935 1.15 0.925 1.27 0.925 1.27 1.165 1.59 1.165 ;
  END
END MXI2X8

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.285 0.29 1.61 ;
        RECT 0.07 1.175 0.22 1.505 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.05 0.815 1.505 ;
        RECT 0.695 1.02 0.815 1.505 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.34 1.515 1.99 ;
        RECT 1.355 0.68 1.475 1.46 ;
        RECT 1.175 0.65 1.435 0.8 ;
        RECT 1.315 0.56 1.435 0.8 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.895 -0.18 1.015 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.625 1.095 2.79 ;
        RECT 0.135 1.745 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.235 1.11 0.935 1.11 0.935 0.9 0.53 0.9 0.53 1.625 0.675 1.625 0.675 1.865 0.555 1.865 0.555 1.745 0.41 1.745 0.41 0.9 0.195 0.9 0.195 0.61 0.315 0.61 0.315 0.78 1.055 0.78 1.055 0.99 1.235 0.99 ;
  END
END AND2X1

MACRO NAND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X2 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.97 2.08 1.09 ;
        RECT 1.84 0.595 1.96 1.09 ;
        RECT 1.81 0.595 1.96 0.855 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.09 ;
        RECT 1.38 1.21 2.84 1.33 ;
        RECT 2.72 0.94 2.84 1.33 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 1.45 3.38 1.57 ;
        RECT 3.26 1.22 3.38 1.57 ;
        RECT 0.96 1.175 1.09 1.57 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.84 1.28 1.09 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 1.69 3.7 1.81 ;
        RECT 3.58 1.22 3.7 1.81 ;
        RECT 3.55 1.465 3.7 1.81 ;
        RECT 0.58 1.22 0.7 1.81 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9696 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.82 1.755 3.99 2.015 ;
        RECT 0.64 1.93 3.94 2.05 ;
        RECT 3.82 0.7 3.94 2.05 ;
        RECT 2.24 0.7 3.94 0.82 ;
        RECT 3.52 1.93 3.64 2.21 ;
        RECT 2.56 1.93 2.68 2.21 ;
        RECT 2.12 0.65 2.36 0.77 ;
        RECT 1.6 1.93 1.72 2.21 ;
        RECT 0.64 1.93 0.76 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.68 0.46 3.92 0.58 ;
        RECT 3.68 -0.18 3.8 0.58 ;
        RECT 0.42 -0.18 0.54 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.94 2.17 4.18 2.29 ;
        RECT 3.94 2.17 4.06 2.79 ;
        RECT 2.98 2.17 3.22 2.29 ;
        RECT 2.98 2.17 3.1 2.79 ;
        RECT 2.02 2.17 2.26 2.29 ;
        RECT 2.02 2.17 2.14 2.79 ;
        RECT 1.06 2.17 1.3 2.29 ;
        RECT 1.06 2.17 1.18 2.79 ;
        RECT 0.22 1.56 0.34 2.79 ;
    END
  END VDD
END NAND4X2

MACRO MX2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 1.255 1.25 1.375 ;
        RECT 0.41 1.695 1.09 1.815 ;
        RECT 0.97 1.255 1.09 1.815 ;
        RECT 0.36 1.475 0.53 1.725 ;
        RECT 0.36 1.465 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.105 0.85 1.575 ;
        RECT 0.73 1.075 0.85 1.575 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.91 1.315 2.25 1.435 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.91 1.315 2.03 1.555 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.175 2.54 1.435 ;
        RECT 2.41 1.175 2.53 2.055 ;
        RECT 2.37 0.475 2.49 1.315 ;
        RECT 2.39 1.175 2.53 1.555 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.89 0.535 2.13 0.655 ;
        RECT 1.89 -0.18 2.01 0.655 ;
        RECT 0.67 -0.18 0.79 0.715 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.99 1.935 2.11 2.79 ;
        RECT 0.71 1.935 0.83 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.25 1.055 1.79 1.055 1.79 1.975 1.53 1.975 1.53 1.995 1.29 1.995 1.29 1.875 1.41 1.875 1.41 1.855 1.67 1.855 1.67 1.055 1.61 1.055 1.61 0.715 1.31 0.715 1.31 0.475 1.43 0.475 1.43 0.595 1.73 0.595 1.73 0.935 2.13 0.935 2.13 0.815 2.25 0.815 ;
      POLYGON 1.55 1.735 1.43 1.735 1.43 1.295 1.37 1.295 1.37 1.075 1.15 1.075 1.15 0.955 0.24 0.955 0.24 1.935 0.41 1.935 0.41 2.175 0.29 2.175 0.29 2.055 0.12 2.055 0.12 0.595 0.25 0.595 0.25 0.475 0.37 0.475 0.37 0.715 0.24 0.715 0.24 0.835 1.49 0.835 1.49 1.175 1.55 1.175 ;
  END
END MX2XL

MACRO TLATNTSCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX3 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.82 0.565 1.09 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.76 1.09 1.18 ;
        RECT 0.925 0.8 1.045 1.24 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.76 1.385 1.24 ;
        RECT 1.23 0.76 1.385 1.215 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.995 0.59 7.115 0.83 ;
        RECT 6.815 0.71 7.115 0.83 ;
        RECT 6.825 1.31 6.945 2.2 ;
        RECT 6.16 0.83 6.935 0.95 ;
        RECT 6.16 1.31 6.945 1.43 ;
        RECT 6.16 0.83 6.31 1.145 ;
        RECT 5.985 1.43 6.28 1.55 ;
        RECT 6.16 0.71 6.28 1.55 ;
        RECT 6.155 0.59 6.275 0.83 ;
        RECT 5.985 1.43 6.105 2.2 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.575 -0.18 6.695 0.64 ;
        RECT 5.675 -0.18 5.795 0.53 ;
        RECT 4.605 -0.18 4.845 0.38 ;
        RECT 3.195 0.7 3.435 0.82 ;
        RECT 3.235 -0.18 3.355 0.82 ;
        RECT 0.985 -0.18 1.105 0.64 ;
        RECT 0.145 -0.18 0.265 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 6.405 1.55 6.525 2.79 ;
        RECT 5.565 1.64 5.685 2.79 ;
        RECT 4.725 1.55 4.845 2.79 ;
        RECT 3.035 2.14 3.275 2.26 ;
        RECT 3.035 2.14 3.155 2.79 ;
        RECT 0.945 1.6 1.065 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.04 1.19 5.565 1.19 5.565 1.52 5.265 1.52 5.265 2.2 5.145 2.2 5.145 1.4 5.445 1.4 5.445 0.92 5.365 0.92 5.365 0.68 5.485 0.68 5.485 0.8 5.565 0.8 5.565 1.07 6.04 1.07 ;
      POLYGON 5.325 1.28 5.125 1.28 5.125 0.62 3.955 0.62 3.955 0.76 3.915 0.76 3.915 1.3 2.955 1.3 2.955 1.66 3.755 1.66 3.755 1.89 3.875 1.89 3.875 2.01 3.635 2.01 3.635 1.78 2.835 1.78 2.835 1.3 2.695 1.3 2.695 1.18 3.795 1.18 3.795 0.64 3.835 0.64 3.835 0.5 5.245 0.5 5.245 1.04 5.325 1.04 ;
      POLYGON 5.005 1.26 4.365 1.26 4.365 1.61 4.485 1.61 4.485 1.73 4.245 1.73 4.245 1.54 3.075 1.54 3.075 1.42 4.245 1.42 4.245 0.86 4.125 0.86 4.125 0.74 4.365 0.74 4.365 1.14 5.005 1.14 ;
      POLYGON 4.585 2.25 3.395 2.25 3.395 2.02 2.515 2.02 2.515 2.07 2.395 2.07 2.395 1.95 2.215 1.95 2.215 0.64 2.335 0.64 2.335 1.83 2.515 1.83 2.515 1.9 3.515 1.9 3.515 2.13 4.465 2.13 4.465 2.01 4.585 2.01 ;
      POLYGON 3.715 0.48 3.675 0.48 3.675 1.06 2.955 1.06 2.955 0.52 2.575 0.52 2.575 1.57 2.715 1.57 2.715 1.69 2.455 1.69 2.455 0.52 1.625 0.52 1.625 1.48 1.545 1.48 1.545 1.72 1.425 1.72 1.425 1.36 1.505 1.36 1.505 0.64 1.405 0.64 1.405 0.4 1.995 0.4 1.995 0.36 2.235 0.36 2.235 0.4 3.075 0.4 3.075 0.94 3.555 0.94 3.555 0.48 3.475 0.48 3.475 0.36 3.715 0.36 ;
      POLYGON 2.095 2.07 1.975 2.07 1.975 1.96 1.185 1.96 1.185 1.48 0.425 1.48 0.425 1.72 0.305 1.72 0.305 1.36 0.685 1.36 0.685 0.7 0.565 0.7 0.565 0.4 0.685 0.4 0.685 0.58 0.805 0.58 0.805 1.36 1.305 1.36 1.305 1.84 1.975 1.84 1.975 0.88 1.795 0.88 1.795 0.64 1.915 0.64 1.915 0.76 2.095 0.76 ;
  END
END TLATNTSCAX3

MACRO AOI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.85 1.67 1.225 ;
        RECT 1.545 0.85 1.665 1.485 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 1.04 0.925 1.295 ;
        RECT 0.65 1.04 0.925 1.16 ;
        RECT 0.65 0.885 0.8 1.16 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.88 2.54 1.35 ;
        RECT 2.39 0.85 2.51 1.35 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.875 0.85 2.085 1.1 ;
        RECT 1.79 0.875 2.025 1.145 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.85 1.38 1.22 ;
        RECT 1.225 1.1 1.345 1.475 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.795 0.51 1.43 ;
        RECT 0.36 0.795 0.51 1.17 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2928 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 1.465 2.83 1.725 ;
        RECT 2.66 0.61 2.78 1.725 ;
        RECT 2.645 1.47 2.765 1.83 ;
        RECT 1.385 0.61 2.78 0.73 ;
        RECT 1.805 1.47 2.83 1.59 ;
        RECT 1.805 1.47 1.925 1.83 ;
        RECT 1.385 0.4 1.505 0.73 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 2.445 0.37 2.685 0.49 ;
        RECT 2.445 -0.18 2.565 0.49 ;
        RECT 0.325 -0.18 0.445 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 0.905 2.23 1.025 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.345 1.95 2.165 1.95 2.165 2.07 1.385 2.07 1.385 1.83 0.485 1.83 0.485 1.71 1.505 1.71 1.505 1.95 2.045 1.95 2.045 1.83 2.225 1.83 2.225 1.71 2.345 1.71 ;
  END
END AOI33XL

MACRO MDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX4 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.185 0.63 2.305 0.87 ;
        RECT 1.965 1.315 2.205 1.65 ;
        RECT 2.085 0.75 2.205 1.65 ;
        RECT 1.23 1.315 2.205 1.435 ;
        RECT 1.345 0.63 1.465 0.87 ;
        RECT 1.005 1.53 1.38 1.65 ;
        RECT 1.23 1.175 1.38 1.65 ;
        RECT 1.26 0.75 1.38 1.65 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.685 1.295 ;
        RECT 0.565 1.055 0.685 1.295 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.595 1.2 7.715 1.44 ;
        RECT 7.32 1.315 7.715 1.435 ;
        RECT 7.32 1.175 7.47 1.435 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.715 1.23 9.06 1.435 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.005 0.99 9.375 1.11 ;
        RECT 8.235 0.97 9.265 1.09 ;
        RECT 9.005 0.94 9.265 1.11 ;
        RECT 8.075 1.19 8.355 1.31 ;
        RECT 8.235 0.97 8.355 1.31 ;
        RECT 8.075 1.19 8.195 1.44 ;
    END
  END S0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.135 -0.18 9.255 0.82 ;
        RECT 7.755 -0.18 7.875 0.83 ;
        RECT 5.465 0.39 5.705 0.51 ;
        RECT 5.585 -0.18 5.705 0.51 ;
        RECT 3.445 -0.18 3.565 0.68 ;
        RECT 2.605 -0.18 2.725 0.68 ;
        RECT 1.765 -0.18 1.885 0.68 ;
        RECT 0.925 -0.18 1.045 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 8.975 1.795 9.095 2.79 ;
        RECT 7.595 1.85 7.715 2.79 ;
        RECT 5.465 2.07 5.705 2.19 ;
        RECT 5.465 2.07 5.585 2.79 ;
        RECT 3.405 2.01 3.645 2.13 ;
        RECT 3.405 2.01 3.525 2.79 ;
        RECT 2.445 2.01 2.685 2.13 ;
        RECT 2.445 2.01 2.565 2.79 ;
        RECT 1.485 2.01 1.725 2.13 ;
        RECT 1.485 2.01 1.605 2.79 ;
        RECT 0.585 2.11 0.705 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.675 0.82 9.615 0.82 9.615 1.68 9.575 1.68 9.575 1.8 9.455 1.8 9.455 1.675 8.475 1.675 8.475 1.24 8.595 1.24 8.595 1.555 9.495 1.555 9.495 0.7 9.555 0.7 9.555 0.58 9.675 0.58 ;
      POLYGON 8.615 0.85 8.115 0.85 8.115 1.07 7.955 1.07 7.955 1.56 8.355 1.56 8.355 2.21 8.235 2.21 8.235 1.68 7.025 1.68 7.025 1.76 6.785 1.76 6.785 1.53 6.905 1.53 6.905 0.72 6.885 0.72 6.885 0.6 7.125 0.6 7.125 0.72 7.025 0.72 7.025 1.56 7.835 1.56 7.835 0.95 7.995 0.95 7.995 0.73 8.495 0.73 8.495 0.59 8.615 0.59 ;
      POLYGON 7.455 0.83 7.335 0.83 7.335 0.48 6.765 0.48 6.765 1.39 6.665 1.39 6.665 1.88 7.235 1.88 7.235 2.03 7.355 2.03 7.355 2.15 7.115 2.15 7.115 2 6.545 2 6.545 1.15 6.645 1.15 6.645 0.48 6.165 0.48 6.165 0.88 6.185 0.88 6.185 1.12 6.045 1.12 6.045 0.75 5.225 0.75 5.225 0.48 4.745 0.48 4.745 1 4.665 1 4.665 1.25 4.125 1.25 4.125 1.37 4.005 1.37 4.005 1.13 4.545 1.13 4.545 0.88 4.625 0.88 4.625 0.36 5.345 0.36 5.345 0.63 6.045 0.63 6.045 0.36 7.455 0.36 ;
      POLYGON 6.525 0.72 6.425 0.72 6.425 1.99 6.305 1.99 6.305 1.36 5.485 1.36 5.485 1.31 5.365 1.31 5.365 1.19 5.605 1.19 5.605 1.24 6.305 1.24 6.305 0.72 6.285 0.72 6.285 0.6 6.525 0.6 ;
      POLYGON 6.265 2.25 6.025 2.25 6.025 1.95 4.925 1.95 4.925 2.23 3.845 2.23 3.845 1.89 0.135 1.89 0.135 1.675 0.12 1.675 0.12 0.935 0.325 0.935 0.325 0.63 0.445 0.63 0.445 1.055 0.24 1.055 0.24 1.555 0.255 1.555 0.255 1.77 3.965 1.77 3.965 2.11 4.805 2.11 4.805 1.23 4.885 1.23 4.885 1.11 5.005 1.11 5.005 1.35 4.925 1.35 4.925 1.83 6.145 1.83 6.145 2.13 6.265 2.13 ;
      POLYGON 5.925 1.07 5.245 1.07 5.245 1.59 5.165 1.59 5.165 1.71 5.045 1.71 5.045 1.47 5.125 1.47 5.125 0.99 4.865 0.99 4.865 0.6 5.105 0.6 5.105 0.87 5.245 0.87 5.245 0.95 5.925 0.95 ;
      POLYGON 4.505 0.72 3.885 0.72 3.885 1.49 4.245 1.49 4.245 1.47 4.365 1.47 4.365 1.99 4.245 1.99 4.245 1.61 3.765 1.61 3.765 1.37 3.185 1.37 3.185 1.13 3.305 1.13 3.305 1.25 3.765 1.25 3.765 0.6 4.505 0.6 ;
      POLYGON 3.645 1.13 3.525 1.13 3.525 1.01 3.065 1.01 3.065 1.53 3.165 1.53 3.165 1.65 2.925 1.65 2.925 1.53 2.945 1.53 2.945 1.01 2.545 1.01 2.545 1.19 2.425 1.19 2.425 0.89 2.945 0.89 2.945 0.66 3.025 0.66 3.025 0.54 3.145 0.54 3.145 0.89 3.645 0.89 ;
  END
END MDFFHQX4

MACRO NOR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.445 0.94 1.815 1.13 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 0.94 2.595 1.09 ;
        RECT 1.215 1.25 2.515 1.37 ;
        RECT 2.395 0.94 2.515 1.37 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 1.49 2.835 1.61 ;
        RECT 2.715 1.22 2.835 1.61 ;
        RECT 0.97 1.28 1.095 1.61 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.855 1.28 1.095 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.02 1.22 3.255 1.46 ;
        RECT 0.495 1.73 3.14 1.85 ;
        RECT 3.02 1.22 3.14 1.85 ;
        RECT 2.97 1.465 3.14 1.85 ;
        RECT 0.495 1.22 0.615 1.85 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.855 1.97 3.495 2.09 ;
        RECT 3.375 0.7 3.495 2.09 ;
        RECT 3.26 1.755 3.495 2.09 ;
        RECT 0.615 0.7 3.495 0.82 ;
        RECT 3.015 0.65 3.255 0.82 ;
        RECT 2.175 0.65 2.415 0.82 ;
        RECT 1.855 1.97 2.095 2.15 ;
        RECT 1.335 0.65 1.575 0.82 ;
        RECT 0.495 0.65 0.735 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.435 0.46 3.675 0.58 ;
        RECT 3.435 -0.18 3.555 0.58 ;
        RECT 2.595 0.46 2.835 0.58 ;
        RECT 2.595 -0.18 2.715 0.58 ;
        RECT 1.755 0.46 1.995 0.58 ;
        RECT 1.755 -0.18 1.875 0.58 ;
        RECT 0.915 0.46 1.155 0.58 ;
        RECT 0.915 -0.18 1.035 0.58 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.195 2.21 3.435 2.79 ;
        RECT 0.435 1.97 0.555 2.79 ;
    END
  END VDD
END NOR4X2

MACRO CLKMX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.605 1.185 1.725 ;
        RECT 1.065 1.31 1.185 1.725 ;
        RECT 0.36 1.465 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 1.28 0.885 1.485 ;
        RECT 0.65 1.09 0.8 1.485 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.905 1.24 2.305 1.38 ;
        RECT 2.045 1.23 2.305 1.38 ;
        RECT 1.905 1.24 2.025 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.175 2.83 1.435 ;
        RECT 2.425 1.175 2.83 1.295 ;
        RECT 2.425 0.59 2.545 1.62 ;
        RECT 2.405 1.5 2.525 2.21 ;
        RECT 2.345 0.47 2.465 0.71 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.765 -0.18 2.885 0.65 ;
        RECT 1.925 -0.18 2.045 0.71 ;
        RECT 0.625 -0.18 0.745 0.71 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.825 1.56 2.945 2.79 ;
        RECT 1.985 1.85 2.105 2.79 ;
        RECT 0.705 1.97 0.825 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.305 1.1 2.065 1.1 2.065 0.95 1.785 0.95 1.785 2.01 1.525 2.01 1.525 2.03 1.285 2.03 1.285 1.91 1.405 1.91 1.405 1.89 1.665 1.89 1.665 0.95 1.425 0.95 1.425 0.73 1.265 0.73 1.265 0.47 1.385 0.47 1.385 0.61 1.545 0.61 1.545 0.83 2.305 0.83 ;
      POLYGON 1.545 1.77 1.425 1.77 1.425 1.19 1.065 1.19 1.065 0.97 0.24 0.97 0.24 1.845 0.405 1.845 0.405 2.09 0.285 2.09 0.285 1.965 0.12 1.965 0.12 0.73 0.205 0.73 0.205 0.47 0.325 0.47 0.325 0.85 1.305 0.85 1.305 1.07 1.545 1.07 ;
  END
END CLKMX2X2

MACRO MX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X6 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 1.555 1.17 1.675 ;
        RECT 1.05 1.35 1.17 1.675 ;
        RECT 0.41 1.195 0.53 1.675 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.045 0.85 1.435 ;
        RECT 0.73 1.035 0.85 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 1.215 2.25 1.435 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.87 1.215 1.99 1.455 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.21 1.43 4.33 2.21 ;
        RECT 3.99 0.8 4.29 0.92 ;
        RECT 4.17 0.405 4.29 0.92 ;
        RECT 4.03 1.43 4.33 1.55 ;
        RECT 4.03 1.19 4.15 1.55 ;
        RECT 3.33 1.04 4.11 1.31 ;
        RECT 3.99 0.8 4.11 1.31 ;
        RECT 3.37 1.04 3.49 2.21 ;
        RECT 3.33 0.405 3.45 1.31 ;
        RECT 2.67 1.19 4.15 1.31 ;
        RECT 2.67 1.175 2.83 1.435 ;
        RECT 2.53 1.36 2.79 1.48 ;
        RECT 2.67 0.63 2.79 1.48 ;
        RECT 2.43 0.63 2.79 0.75 ;
        RECT 2.53 1.36 2.65 2.21 ;
        RECT 2.43 0.4 2.55 0.75 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.75 -0.18 3.87 0.92 ;
        RECT 2.91 -0.18 3.03 0.92 ;
        RECT 2.01 -0.18 2.13 0.74 ;
        RECT 0.73 -0.18 0.85 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.79 1.43 3.91 2.79 ;
        RECT 2.95 1.43 3.07 2.79 ;
        RECT 2.11 1.555 2.23 2.79 ;
        RECT 0.57 1.795 0.69 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.49 1.24 2.37 1.24 2.37 0.99 1.75 0.99 1.75 1.84 1.43 1.84 1.43 2.21 1.31 2.21 1.31 1.72 1.63 1.72 1.63 0.99 1.47 0.99 1.47 0.675 1.37 0.675 1.37 0.435 1.49 0.435 1.49 0.555 1.59 0.555 1.59 0.87 2.49 0.87 ;
      POLYGON 1.51 1.6 1.39 1.6 1.39 1.23 1.23 1.23 1.23 0.915 0.24 0.915 0.24 1.555 0.27 1.555 0.27 2.035 0.15 2.035 0.15 1.675 0.12 1.675 0.12 0.675 0.25 0.675 0.25 0.5 0.37 0.5 0.37 0.795 1.35 0.795 1.35 1.11 1.51 1.11 ;
  END
END MX2X6

MACRO MXI2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X6 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 1.555 1.19 1.675 ;
        RECT 1.07 1.095 1.19 1.675 ;
        RECT 0.41 1.315 0.53 1.675 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.095 0.87 1.42 ;
        RECT 0.65 1.105 0.835 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.89 1.175 2.25 1.415 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.03 0.405 5.15 1.04 ;
        RECT 4.95 1.19 5.07 2.21 ;
        RECT 4.85 0.92 5.15 1.04 ;
        RECT 4.19 1.04 4.97 1.31 ;
        RECT 4.19 0.405 4.31 1.31 ;
        RECT 4.11 1.19 4.23 2.21 ;
        RECT 3.55 1.19 5.07 1.31 ;
        RECT 3.55 1.175 3.7 1.435 ;
        RECT 3.29 1.07 3.67 1.19 ;
        RECT 3.27 1.31 3.7 1.43 ;
        RECT 3.29 0.4 3.41 1.19 ;
        RECT 3.27 1.31 3.39 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.61 -0.18 4.73 0.92 ;
        RECT 3.77 -0.18 3.89 0.92 ;
        RECT 2.87 -0.18 2.99 0.845 ;
        RECT 2.03 -0.18 2.15 0.655 ;
        RECT 0.75 -0.18 0.87 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.53 1.43 4.65 2.79 ;
        RECT 3.69 1.555 3.81 2.79 ;
        RECT 2.85 1.56 2.97 2.79 ;
        RECT 2.01 1.675 2.13 2.79 ;
        RECT 0.67 1.795 0.79 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.15 1.26 2.73 1.26 2.73 1.68 2.55 1.68 2.55 2.21 2.43 2.21 2.43 1.56 2.61 1.56 2.61 0.815 2.45 0.815 2.45 0.575 2.57 0.575 2.57 0.695 2.73 0.695 2.73 1.14 3.15 1.14 ;
      POLYGON 2.49 1.175 2.37 1.175 2.37 1.055 1.77 1.055 1.77 1.815 1.49 1.815 1.49 1.915 1.25 1.915 1.25 1.795 1.37 1.795 1.37 1.695 1.65 1.695 1.65 1.055 1.55 1.055 1.55 0.655 1.39 0.655 1.39 0.415 1.51 0.415 1.51 0.535 1.67 0.535 1.67 0.935 2.49 0.935 ;
      POLYGON 1.53 1.575 1.41 1.575 1.41 1.295 1.31 1.295 1.31 0.975 0.24 0.975 0.24 1.555 0.29 1.555 0.29 1.915 0.17 1.915 0.17 1.675 0.12 1.675 0.12 0.535 0.33 0.535 0.33 0.415 0.45 0.415 0.45 0.655 0.24 0.655 0.24 0.855 1.31 0.855 1.31 0.775 1.43 0.775 1.43 1.175 1.53 1.175 ;
  END
END MXI2X6

MACRO BUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.685 1.26 7.285 1.38 ;
        RECT 6.685 1.23 6.945 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.565 0.715 5.805 0.835 ;
        RECT 5.625 1.295 5.745 2.21 ;
        RECT 0.545 0.765 5.685 0.885 ;
        RECT 0.545 1.295 5.745 1.415 ;
        RECT 4.725 0.715 4.965 0.885 ;
        RECT 4.785 1.295 4.905 2.21 ;
        RECT 3.885 0.715 4.125 0.885 ;
        RECT 3.945 1.295 4.065 2.21 ;
        RECT 3.045 0.715 3.285 0.885 ;
        RECT 3.105 1.295 3.225 2.21 ;
        RECT 2.205 0.715 2.445 0.885 ;
        RECT 2.265 1.295 2.385 2.21 ;
        RECT 1.365 0.715 1.605 0.885 ;
        RECT 1.425 1.295 1.545 2.21 ;
        RECT 0.585 1.295 0.8 1.725 ;
        RECT 0.585 1.295 0.705 2.21 ;
        RECT 0.585 0.645 0.705 0.885 ;
        RECT 0.545 0.765 0.665 1.415 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.725 -0.18 7.845 0.705 ;
        RECT 6.885 -0.18 7.005 0.705 ;
        RECT 6.045 -0.18 6.165 0.705 ;
        RECT 5.205 -0.18 5.325 0.645 ;
        RECT 4.365 -0.18 4.485 0.645 ;
        RECT 3.525 -0.18 3.645 0.645 ;
        RECT 2.685 -0.18 2.805 0.645 ;
        RECT 1.845 -0.18 1.965 0.645 ;
        RECT 1.005 -0.18 1.125 0.64 ;
        RECT 0.165 -0.18 0.285 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.725 1.56 7.845 2.79 ;
        RECT 6.885 1.74 7.005 2.79 ;
        RECT 6.045 1.56 6.165 2.79 ;
        RECT 5.205 1.535 5.325 2.79 ;
        RECT 4.365 1.535 4.485 2.79 ;
        RECT 3.525 1.535 3.645 2.79 ;
        RECT 2.685 1.535 2.805 2.79 ;
        RECT 1.845 1.535 1.965 2.79 ;
        RECT 1.005 1.535 1.125 2.79 ;
        RECT 0.165 1.465 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.425 0.945 6.565 0.945 6.565 1.5 7.425 1.5 7.425 2.21 7.305 2.21 7.305 1.62 6.585 1.62 6.585 2.21 6.465 2.21 6.465 1.62 6.445 1.62 6.445 1.175 0.785 1.175 0.785 1.055 6.445 1.055 6.445 0.825 6.465 0.825 6.465 0.655 6.585 0.655 6.585 0.825 7.305 0.825 7.305 0.655 7.425 0.655 ;
  END
END BUFX16

MACRO XOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X1 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4014 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.27 1.56 8.51 2.25 ;
        RECT 8.39 0.36 8.51 2.25 ;
        RECT 8.135 0.65 8.51 0.8 ;
        RECT 8.27 0.36 8.51 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.099 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.07 0.325 1.47 ;
        RECT 0.07 1.175 0.325 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3198 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.267 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.1978 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.23 1.145 1.38 ;
        RECT 0.845 1.03 1.025 1.375 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 1.35 6.81 1.47 ;
        RECT 6.08 1.23 6.365 1.47 ;
        RECT 6.08 0.905 6.2 1.47 ;
        RECT 5.695 0.905 6.2 1.025 ;
    END
  END C
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.73 2.29 7.97 2.79 ;
        RECT 7.79 1.69 7.91 2.79 ;
        RECT 1.865 2.27 2.105 2.79 ;
        RECT 0.685 2.29 0.925 2.79 ;
        RECT 0.745 1.97 0.865 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.73 -0.18 7.97 0.32 ;
        RECT 7.79 -0.18 7.91 0.67 ;
        RECT 1.865 -0.18 2.105 0.32 ;
        RECT 0.685 -0.18 0.925 0.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.23 1.315 7.67 1.315 7.67 2.17 6.26 2.17 6.26 1.89 6.56 1.89 6.56 2.05 7.55 2.05 7.55 0.62 7.42 0.62 7.42 0.48 6.26 0.48 6.26 0.36 7.54 0.36 7.54 0.5 7.67 0.5 7.67 1.195 7.99 1.195 7.99 1.075 8.23 1.075 ;
      POLYGON 7.43 0.86 7.345 0.86 7.345 1.81 7.43 1.81 7.43 1.93 7.19 1.93 7.19 1.81 7.225 1.81 7.225 0.86 7.19 0.86 7.19 0.74 7.43 0.74 ;
      POLYGON 7.05 1.77 7.04 1.77 7.04 1.79 6.8 1.79 6.8 1.77 4.275 1.77 4.275 1.65 5.095 1.65 5.095 0.72 4.525 0.72 4.525 0.6 5.215 0.6 5.215 1.65 6.93 1.65 6.93 0.72 6.8 0.72 6.8 0.6 7.05 0.6 ;
      POLYGON 5.96 0.705 5.9 0.705 5.9 0.72 5.48 0.72 5.48 1.405 5.96 1.405 5.96 1.525 5.36 1.525 5.36 0.6 5.72 0.6 5.72 0.585 5.96 0.585 ;
      RECT 2.985 1.89 5.96 2.01 ;
      RECT 2.405 0.36 5.64 0.48 ;
      RECT 2.405 2.13 5.64 2.25 ;
      POLYGON 4.97 1.04 4.17 1.04 4.17 1.285 4.05 1.285 4.05 0.92 4.97 0.92 ;
      POLYGON 4.075 0.72 3.93 0.72 3.93 1.77 1.725 1.77 1.725 2.17 0.985 2.17 0.985 1.81 0.325 1.81 0.325 1.93 0.205 1.93 0.205 1.69 0.505 1.69 0.505 0.92 0.205 0.92 0.205 0.44 1.605 0.44 1.605 0.32 1.725 0.32 1.725 0.56 0.325 0.56 0.325 0.8 0.625 0.8 0.625 1.69 1.105 1.69 1.105 2.05 1.605 2.05 1.605 1.65 3.81 1.65 3.81 0.6 4.075 0.6 ;
      POLYGON 3.69 1.08 3.57 1.08 3.57 1.02 2.81 1.02 2.81 1.16 2.885 1.16 2.885 1.28 2.645 1.28 2.645 1.16 2.69 1.16 2.69 0.9 3.57 0.9 3.57 0.84 3.69 0.84 ;
      POLYGON 3.225 1.53 1.94 1.53 1.94 0.6 3.205 0.6 3.205 0.72 2.06 0.72 2.06 1.41 3.225 1.41 ;
      POLYGON 1.485 1.12 1.405 1.12 1.405 1.81 1.465 1.81 1.465 1.93 1.225 1.93 1.225 1.81 1.285 1.81 1.285 1.12 1.245 1.12 1.245 1 1.285 1 1.285 0.8 1.225 0.8 1.225 0.68 1.465 0.68 1.465 0.8 1.405 0.8 1.405 1 1.485 1 ;
  END
END XOR3X1

MACRO TLATSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRXL 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 1.255 2.305 1.475 ;
        RECT 2.045 1.23 2.305 1.475 ;
    END
  END SN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.765 1.27 2.885 1.595 ;
        RECT 2.68 1.455 2.83 1.725 ;
    END
  END G
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.15 4.045 1.41 ;
        RECT 3.765 1.15 4.045 1.39 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 1.465 5.915 1.61 ;
        RECT 5.795 1.26 5.915 1.61 ;
        RECT 5.58 1.465 5.73 1.815 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 1.83 ;
        RECT 1.23 1.465 1.485 1.725 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 5.955 -0.18 6.075 0.78 ;
        RECT 3.985 0.43 4.225 0.55 ;
        RECT 4.105 -0.18 4.225 0.55 ;
        RECT 1.725 0.74 1.965 0.86 ;
        RECT 1.725 -0.18 1.845 0.86 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 5.875 2.2 6.115 2.79 ;
        RECT 4.365 2.01 4.485 2.79 ;
        RECT 3.525 2.23 3.645 2.79 ;
        RECT 2.685 2.23 2.805 2.79 ;
        RECT 1.845 2.23 1.965 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.535 1.84 6.415 1.84 6.415 1.72 6.375 1.72 6.375 1.14 5.595 1.14 5.595 1.2 5.475 1.2 5.475 0.96 5.595 0.96 5.595 1.02 6.375 1.02 6.375 0.54 6.495 0.54 6.495 1.6 6.535 1.6 ;
      POLYGON 6.475 2.22 6.235 2.22 6.235 2.08 5.555 2.08 5.555 2.22 5.315 2.22 5.315 2.08 4.995 2.08 4.995 1.04 4.875 1.04 4.875 1.03 3.465 1.03 3.465 1.71 3.165 1.71 3.165 1.83 3.045 1.83 3.045 1.59 3.345 1.59 3.345 0.72 3.285 0.72 3.285 0.6 3.525 0.6 3.525 0.72 3.465 0.72 3.465 0.91 5.115 0.91 5.115 1.96 6.355 1.96 6.355 2.1 6.475 2.1 ;
      POLYGON 5.355 1.84 5.235 1.84 5.235 0.79 3.67 0.79 3.67 0.48 2.995 0.48 2.995 0.54 2.225 0.54 2.225 0.42 2.875 0.42 2.875 0.36 3.79 0.36 3.79 0.67 5.215 0.67 5.215 0.54 5.335 0.54 5.335 0.66 5.355 0.66 ;
      POLYGON 4.875 1.8 4.755 1.8 4.755 1.89 3.825 1.89 3.825 1.77 4.635 1.77 4.635 1.68 4.875 1.68 ;
      POLYGON 4.285 1.65 3.705 1.65 3.705 2.07 2.735 2.07 2.735 1.965 2.205 1.965 2.205 1.605 2.425 1.605 2.425 1.11 1.745 1.11 1.745 1.26 1.625 1.26 1.625 0.99 2.425 0.99 2.425 0.68 2.545 0.68 2.545 1.725 2.325 1.725 2.325 1.845 2.855 1.845 2.855 1.95 3.585 1.95 3.585 1.53 4.165 1.53 4.165 1.27 4.285 1.27 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END TLATSRXL

MACRO OAI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X1 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.28 1.3 1.52 1.42 ;
        RECT 1.28 0.595 1.4 1.42 ;
        RECT 1.23 0.595 1.4 0.855 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 1.195 1.16 1.4 ;
        RECT 0.94 1.04 1.09 1.435 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.04 0.8 1.435 ;
        RECT 0.56 1.115 0.8 1.32 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.4 1.4 ;
        RECT 0.28 1.16 0.4 1.4 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5104 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.555 1.76 1.675 ;
        RECT 1.64 0.75 1.76 1.675 ;
        RECT 1.62 1.555 1.74 2.21 ;
        RECT 1.62 0.63 1.74 0.87 ;
        RECT 1.52 1.555 1.74 2.015 ;
        RECT 0.78 1.555 0.9 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 0.56 -0.18 0.68 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.2 1.795 1.32 2.79 ;
        RECT 0.14 1.56 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.1 0.92 0.14 0.92 0.14 0.63 0.26 0.63 0.26 0.8 0.98 0.8 0.98 0.63 1.1 0.63 ;
  END
END OAI211X1

MACRO TBUFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFXL 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 1.16 1.415 1.28 ;
        RECT 0.435 1.025 0.8 1.28 ;
        RECT 0.65 0.885 0.8 1.28 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.22 0.36 2.725 0.48 ;
        RECT 1.215 0.44 2.34 0.56 ;
        RECT 0.815 1.4 1.655 1.52 ;
        RECT 1.535 0.92 1.655 1.52 ;
        RECT 1.215 0.92 1.655 1.04 ;
        RECT 1.175 1.4 1.435 1.67 ;
        RECT 1.215 0.44 1.335 1.04 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.245 0.76 3.365 1.605 ;
        RECT 2.97 1.465 3.345 1.725 ;
        RECT 3.225 0.64 3.345 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.845 -0.18 2.965 0.76 ;
        RECT 2.805 0.64 2.925 0.88 ;
        RECT 1.845 -0.18 2.085 0.32 ;
        RECT 0.975 -0.18 1.095 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.745 2.085 2.865 2.79 ;
        RECT 1.035 2.29 1.275 2.79 ;
        RECT 0.135 1.88 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.185 2.185 3.065 2.185 3.065 1.965 2.39 1.965 2.39 2.17 1.21 2.17 1.21 2.11 0.615 2.11 0.615 1.76 0.195 1.76 0.195 0.785 0.275 0.785 0.275 0.62 0.395 0.62 0.395 0.905 0.315 0.905 0.315 1.64 0.735 1.64 0.735 1.99 1.33 1.99 1.33 2.05 2.27 2.05 2.27 1.845 3.185 1.845 ;
      POLYGON 3.125 1.14 2.525 1.14 2.525 1.485 2.165 1.485 2.165 1.725 2.045 1.725 2.045 1.365 2.405 1.365 2.405 0.82 2.325 0.82 2.325 0.7 2.565 0.7 2.565 0.82 2.525 0.82 2.525 1.02 3.125 1.02 ;
      POLYGON 2.285 1.245 1.895 1.245 1.895 1.93 1.515 1.93 1.515 1.81 1.775 1.81 1.775 0.8 1.455 0.8 1.455 0.68 1.895 0.68 1.895 1.125 2.285 1.125 ;
  END
END TBUFXL

MACRO DFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 0.92 7.525 1.19 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.255 2.105 1.46 ;
        RECT 1.755 1.23 2.015 1.46 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3312 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.76 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.195 3.275 1.395 ;
        RECT 2.915 1.17 3.175 1.395 ;
    END
  END RN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2888 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.375 0.61 1.495 0.87 ;
        RECT 1.285 1.23 1.405 2.21 ;
        RECT 1.265 0.75 1.385 1.35 ;
        RECT 1.23 0.885 1.385 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.265 0.68 7.505 0.8 ;
        RECT 7.385 -0.18 7.505 0.8 ;
        RECT 5.425 0.47 5.665 0.59 ;
        RECT 5.545 -0.18 5.665 0.59 ;
        RECT 3.315 0.61 3.555 0.73 ;
        RECT 3.435 -0.18 3.555 0.73 ;
        RECT 1.735 0.67 1.975 0.79 ;
        RECT 1.735 -0.18 1.855 0.79 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.665 2.11 7.785 2.79 ;
        RECT 6.065 2.15 6.185 2.79 ;
        RECT 5.255 2.29 5.495 2.79 ;
        RECT 3.375 2.29 3.615 2.79 ;
        RECT 2.515 2.15 2.635 2.79 ;
        RECT 1.765 2.2 1.885 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.325 1.75 8.085 1.75 8.085 1.43 7.225 1.43 7.225 1.55 7.105 1.55 7.105 1.43 7.025 1.43 7.025 0.5 5.905 0.5 5.905 0.83 5.185 0.83 5.185 0.49 4.705 0.49 4.705 1.07 4.055 1.07 4.055 1.41 3.935 1.41 3.935 0.95 4.585 0.95 4.585 0.37 5.305 0.37 5.305 0.71 5.785 0.71 5.785 0.38 6.235 0.38 6.235 0.36 6.475 0.36 6.475 0.38 7.145 0.38 7.145 1.31 7.825 1.31 7.825 0.62 7.945 0.62 7.945 1.31 8.205 1.31 8.205 1.63 8.325 1.63 ;
      POLYGON 8.125 2.25 8.005 2.25 8.005 1.99 7.33 1.99 7.33 2.15 6.92 2.15 6.92 2.25 6.68 2.25 6.68 2.15 6.305 2.15 6.305 1.93 2.125 1.93 2.125 1.58 2.335 1.58 2.335 0.61 2.455 0.61 2.455 1.81 4.595 1.81 4.595 1.31 4.815 1.31 4.815 1.19 4.935 1.19 4.935 1.43 4.715 1.43 4.715 1.81 6.425 1.81 6.425 2.03 7.21 2.03 7.21 1.87 8.125 1.87 ;
      POLYGON 7.085 1.91 6.965 1.91 6.965 1.79 6.865 1.79 6.865 1.67 6.785 1.67 6.785 1.36 5.415 1.36 5.415 1.43 5.295 1.43 5.295 1.19 5.415 1.19 5.415 1.24 6.545 1.24 6.545 0.62 6.665 0.62 6.665 1.24 6.905 1.24 6.905 1.55 6.985 1.55 6.985 1.67 7.085 1.67 ;
      POLYGON 6.665 1.87 6.545 1.87 6.545 1.69 5.735 1.69 5.735 1.57 6.665 1.57 ;
      POLYGON 6.225 1.12 5.985 1.12 5.985 1.07 5.175 1.07 5.175 1.69 4.835 1.69 4.835 1.57 5.055 1.57 5.055 1.07 4.825 1.07 4.825 0.61 5.065 0.61 5.065 0.95 6.105 0.95 6.105 1 6.225 1 ;
      RECT 3.055 2.05 5.815 2.17 ;
      POLYGON 4.465 0.73 3.815 0.73 3.815 1.53 4.155 1.53 4.155 1.57 4.275 1.57 4.275 1.69 4.035 1.69 4.035 1.65 3.695 1.65 3.695 1.05 2.815 1.05 2.815 0.93 3.695 0.93 3.695 0.61 4.465 0.61 ;
      POLYGON 3.575 1.635 3.135 1.635 3.135 1.69 2.895 1.69 2.895 1.635 2.575 1.635 2.575 0.67 2.735 0.67 2.735 0.49 2.215 0.49 2.215 1.11 1.505 1.11 1.505 0.99 2.095 0.99 2.095 0.37 2.855 0.37 2.855 0.79 2.695 0.79 2.695 1.515 3.455 1.515 3.455 1.19 3.575 1.19 ;
      POLYGON 1.105 0.92 1.095 0.92 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.8 0.985 0.8 0.985 0.68 1.105 0.68 ;
  END
END DFFRX1

MACRO AND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.06 0.24 1.515 ;
        RECT 0.12 1.04 0.24 1.515 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.04 0.87 1.35 ;
        RECT 0.36 1.12 0.87 1.24 ;
        RECT 0.36 1.12 0.51 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.12 1.38 1.575 ;
        RECT 1.23 1.09 1.35 1.575 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.93 1.145 2.05 2.01 ;
        RECT 1.81 0.885 1.96 1.265 ;
        RECT 1.81 0.68 1.93 1.265 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.39 -0.18 1.51 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.51 1.575 1.63 2.79 ;
        RECT 0.615 2.215 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 1.26 1.57 1.26 1.57 0.97 1.11 0.97 1.11 1.695 1.21 1.695 1.21 1.935 1.09 1.935 1.09 1.815 0.99 1.815 0.99 1.755 0.075 1.755 0.075 1.635 0.99 1.635 0.99 0.92 0.27 0.92 0.27 0.68 0.39 0.68 0.39 0.8 1.11 0.8 1.11 0.85 1.69 0.85 ;
  END
END AND3X1

MACRO OAI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X2 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.15 1.155 3.465 1.38 ;
        RECT 2.97 1.155 3.465 1.355 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.505 1.01 4.625 1.42 ;
        RECT 4.365 1.15 4.625 1.38 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.165 1.215 1.38 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.225 5.445 1.345 ;
        RECT 5 1.175 5.15 1.435 ;
        RECT 4.085 1.54 5.12 1.66 ;
        RECT 5 1.175 5.12 1.66 ;
        RECT 4.085 1.22 4.205 1.66 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.5 3.785 1.62 ;
        RECT 3.665 1.22 3.785 1.62 ;
        RECT 2.68 1.175 2.83 1.62 ;
        RECT 2.445 1.28 2.83 1.4 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.535 1.5 1.715 1.62 ;
        RECT 1.52 1.22 1.715 1.62 ;
        RECT 1.52 1.175 1.67 1.62 ;
        RECT 0.535 1.22 0.655 1.62 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.565 1.465 5.73 1.725 ;
        RECT 1.115 1.78 5.685 1.9 ;
        RECT 5.565 0.77 5.685 1.9 ;
        RECT 4.345 0.77 5.685 0.89 ;
        RECT 5.185 0.6 5.305 0.89 ;
        RECT 4.565 1.78 4.685 2.21 ;
        RECT 4.345 0.6 4.465 0.89 ;
        RECT 2.985 1.74 3.105 2.21 ;
        RECT 1.115 1.74 1.235 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 1.855 -0.18 1.975 0.73 ;
        RECT 1.015 -0.18 1.135 0.73 ;
        RECT 0.175 -0.18 0.295 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.145 2.02 5.385 2.15 ;
        RECT 5.145 2.02 5.265 2.79 ;
        RECT 3.865 2.02 4.105 2.15 ;
        RECT 3.865 2.02 3.985 2.79 ;
        RECT 2.185 2.02 2.425 2.15 ;
        RECT 2.185 2.02 2.305 2.79 ;
        RECT 0.375 1.74 0.495 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.725 0.65 5.605 0.65 5.605 0.48 4.885 0.48 4.885 0.65 4.765 0.65 4.765 0.48 4.045 0.48 4.045 0.65 3.925 0.65 3.925 0.48 3.205 0.48 3.205 0.65 3.085 0.65 3.085 0.48 2.365 0.48 2.365 0.65 2.245 0.65 2.245 0.36 5.725 0.36 ;
      POLYGON 3.625 0.97 0.595 0.97 0.595 0.68 0.715 0.68 0.715 0.85 1.435 0.85 1.435 0.68 1.555 0.68 1.555 0.85 2.665 0.85 2.665 0.6 2.785 0.6 2.785 0.85 3.505 0.85 3.505 0.6 3.625 0.6 ;
  END
END OAI222X2

MACRO OAI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X4 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.26 8.855 1.38 ;
        RECT 7.845 1.23 8.105 1.38 ;
        RECT 7.955 1 8.075 1.38 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.435 ;
        RECT 1.535 0.94 1.655 1.435 ;
        RECT 0.895 1.28 1.67 1.4 ;
        RECT 0.775 1.3 1.015 1.42 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.535 1.22 5.095 1.34 ;
        RECT 4.655 1.22 4.915 1.38 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.175 3.41 1.435 ;
        RECT 3.26 0.94 3.38 1.435 ;
        RECT 2.435 1.28 3.41 1.4 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.215 1.22 6.775 1.34 ;
        RECT 6.395 1.22 6.655 1.38 ;
    END
  END B2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.655 1.26 10.555 1.38 ;
        RECT 9.655 1.23 10.135 1.38 ;
        RECT 9.655 1 9.775 1.38 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.8136 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.155 0.65 10.395 0.77 ;
        RECT 5.955 0.76 10.275 0.88 ;
        RECT 9.315 0.65 9.555 0.88 ;
        RECT 8.475 0.65 8.715 0.88 ;
        RECT 7.635 0.65 7.875 0.88 ;
        RECT 7.275 1.5 7.395 2.01 ;
        RECT 3.915 1.5 7.395 1.62 ;
        RECT 6.795 0.65 7.035 0.88 ;
        RECT 6.435 1.5 6.555 2.01 ;
        RECT 5.955 0.65 6.195 0.88 ;
        RECT 4.215 0.98 6.075 1.1 ;
        RECT 5.955 0.65 6.075 1.1 ;
        RECT 5.595 1.5 5.715 2.15 ;
        RECT 4.755 1.5 4.875 2.01 ;
        RECT 4.215 0.98 4.335 1.62 ;
        RECT 4.075 1.23 4.335 1.38 ;
        RECT 3.915 1.5 4.035 2.01 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 5.115 0.46 5.355 0.58 ;
        RECT 5.115 -0.18 5.235 0.58 ;
        RECT 4.275 0.46 4.515 0.58 ;
        RECT 4.275 -0.18 4.395 0.58 ;
        RECT 3.435 0.46 3.675 0.58 ;
        RECT 3.435 -0.18 3.555 0.58 ;
        RECT 2.595 0.46 2.835 0.58 ;
        RECT 2.595 -0.18 2.715 0.58 ;
        RECT 1.755 0.46 1.995 0.58 ;
        RECT 1.755 -0.18 1.875 0.58 ;
        RECT 0.915 0.46 1.155 0.58 ;
        RECT 0.915 -0.18 1.035 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.635 1.74 10.755 2.79 ;
        RECT 9.795 1.74 9.915 2.79 ;
        RECT 1.395 1.795 1.515 2.79 ;
        RECT 0.555 1.795 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.175 2.21 11.055 2.21 11.055 1.62 10.335 1.62 10.335 2.21 10.215 2.21 10.215 1.62 9.495 1.62 9.495 2.21 9.375 2.21 9.375 1.62 8.655 1.62 8.655 2.01 8.535 2.01 8.535 1.62 7.815 1.62 7.815 2.01 7.695 2.01 7.695 1.5 11.175 1.5 ;
      POLYGON 10.755 0.65 10.635 0.65 10.635 0.53 9.915 0.53 9.915 0.64 9.795 0.64 9.795 0.53 9.075 0.53 9.075 0.64 8.955 0.64 8.955 0.53 8.235 0.53 8.235 0.64 8.115 0.64 8.115 0.53 7.395 0.53 7.395 0.64 7.275 0.64 7.275 0.53 6.555 0.53 6.555 0.64 6.435 0.64 6.435 0.53 5.715 0.53 5.715 0.82 0.555 0.82 0.555 0.58 0.675 0.58 0.675 0.7 1.395 0.7 1.395 0.58 1.515 0.58 1.515 0.7 2.235 0.7 2.235 0.58 2.355 0.58 2.355 0.7 3.075 0.7 3.075 0.58 3.195 0.58 3.195 0.7 3.915 0.7 3.915 0.58 4.035 0.58 4.035 0.7 4.755 0.7 4.755 0.58 4.875 0.58 4.875 0.7 5.595 0.7 5.595 0.41 6.435 0.41 6.435 0.4 6.555 0.4 6.555 0.41 7.275 0.41 7.275 0.4 7.395 0.4 7.395 0.41 8.115 0.41 8.115 0.4 8.235 0.4 8.235 0.41 8.955 0.41 8.955 0.4 9.075 0.4 9.075 0.41 9.795 0.41 9.795 0.4 9.915 0.4 9.915 0.41 10.755 0.41 ;
      POLYGON 9.075 2.25 6.015 2.25 6.015 1.74 6.135 1.74 6.135 2.13 6.855 2.13 6.855 1.74 6.975 1.74 6.975 2.13 8.115 2.13 8.115 1.74 8.235 1.74 8.235 2.13 8.955 2.13 8.955 1.74 9.075 1.74 ;
      POLYGON 5.295 2.25 2.235 2.25 2.235 1.795 2.355 1.795 2.355 2.13 3.075 2.13 3.075 1.795 3.195 1.795 3.195 2.13 4.335 2.13 4.335 1.74 4.455 1.74 4.455 2.13 5.175 2.13 5.175 1.74 5.295 1.74 ;
      POLYGON 3.615 2.01 3.495 2.01 3.495 1.675 2.775 1.675 2.775 2.01 2.655 2.01 2.655 1.675 1.935 1.675 1.935 2.21 1.815 2.21 1.815 1.675 1.095 1.675 1.095 2.21 0.975 2.21 0.975 1.675 0.255 1.675 0.255 2.21 0.135 2.21 0.135 1.555 3.615 1.555 ;
  END
END OAI33X4

MACRO MXI2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X4 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.595 0.935 1.715 1.755 ;
        RECT 0.955 1.635 1.715 1.755 ;
        RECT 1.035 1.505 1.155 1.755 ;
        RECT 0.39 1.725 1.075 1.845 ;
        RECT 0.36 1.465 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.175 0.835 1.605 ;
        RECT 0.65 1.175 0.835 1.59 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.075 1.05 2.25 1.48 ;
        RECT 2.075 1.03 2.195 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.635 0.68 3.835 0.8 ;
        RECT 3.455 1.32 3.575 2.21 ;
        RECT 2.625 1.32 3.575 1.44 ;
        RECT 2.625 1.23 2.885 1.44 ;
        RECT 2.615 1.44 2.875 1.56 ;
        RECT 2.755 0.68 2.875 1.56 ;
        RECT 2.615 1.44 2.735 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.195 0.49 4.435 0.61 ;
        RECT 4.315 -0.18 4.435 0.61 ;
        RECT 3.115 -0.18 3.355 0.32 ;
        RECT 2.155 -0.18 2.275 0.67 ;
        RECT 0.655 -0.18 0.775 0.815 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 3.875 1.56 3.995 2.79 ;
        RECT 3.035 1.56 3.155 2.79 ;
        RECT 2.195 1.6 2.315 2.79 ;
        RECT 0.555 1.965 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.795 0.86 4.515 0.86 4.515 1.42 4.415 1.42 4.415 2.21 4.295 2.21 4.295 1.42 3.695 1.42 3.695 1.3 4.395 1.3 4.395 0.74 4.675 0.74 4.675 0.62 4.795 0.62 ;
      POLYGON 4.275 1.18 4.155 1.18 4.155 0.85 3.955 0.85 3.955 0.56 2.515 0.56 2.515 0.91 1.955 0.91 1.955 2.085 1.315 2.085 1.315 2.205 1.195 2.205 1.195 1.965 1.835 1.965 1.835 0.815 1.455 0.815 1.455 0.575 1.575 0.575 1.575 0.695 1.955 0.695 1.955 0.79 2.395 0.79 2.395 0.44 4.075 0.44 4.075 0.73 4.275 0.73 ;
      POLYGON 1.475 1.515 1.355 1.515 1.355 1.055 0.24 1.055 0.24 1.845 0.255 1.845 0.255 2.085 0.135 2.085 0.135 1.965 0.12 1.965 0.12 0.815 0.235 0.815 0.235 0.575 0.355 0.575 0.355 0.935 1.475 0.935 ;
  END
END MXI2X4

MACRO CLKAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.151 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.04 1.59 1.16 ;
        RECT 0.595 0.99 1.385 1.11 ;
        RECT 0.595 0.94 0.855 1.11 ;
        RECT 0.39 1.04 0.715 1.16 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.151 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 1.255 1.145 1.48 ;
        RECT 0.885 1.23 1.145 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.03 1.29 3.15 2.18 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 2.97 0.76 3.09 1.435 ;
        RECT 2.19 1.29 3.15 1.41 ;
        RECT 1.99 0.81 3.09 0.93 ;
        RECT 2.83 0.76 3.09 0.93 ;
        RECT 2.83 0.64 2.95 0.93 ;
        RECT 2.19 1.29 2.31 2.18 ;
        RECT 1.99 0.64 2.11 0.93 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.25 -0.18 3.37 0.69 ;
        RECT 2.41 -0.18 2.53 0.69 ;
        RECT 1.51 0.51 1.75 0.63 ;
        RECT 1.51 -0.18 1.63 0.63 ;
        RECT 0.29 -0.18 0.41 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.45 1.53 3.57 2.79 ;
        RECT 2.61 1.53 2.73 2.79 ;
        RECT 1.71 2.135 1.83 2.79 ;
        RECT 0.87 2.135 0.99 2.79 ;
        RECT 0.135 2.135 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.85 1.17 1.83 1.17 1.83 1.72 0.45 1.72 0.45 1.6 1.71 1.6 1.71 0.87 0.99 0.87 0.99 0.82 0.87 0.82 0.87 0.7 1.11 0.7 1.11 0.75 1.83 0.75 1.83 1.05 2.85 1.05 ;
  END
END CLKAND2X4

MACRO DFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX1 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.135 1.2 3.465 1.415 ;
        RECT 3.015 1.2 3.465 1.39 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.035 1.22 8.155 1.51 ;
        RECT 7.9 1.175 8.05 1.475 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 1.04 8.63 1.435 ;
        RECT 8.495 0.835 8.615 1.435 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.66 1.485 1.99 ;
        RECT 1.23 0.885 1.485 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.375 -0.18 8.495 0.38 ;
        RECT 6.605 -0.18 6.845 0.32 ;
        RECT 3.295 -0.18 3.415 0.38 ;
        RECT 1.845 -0.18 1.965 0.38 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.195 1.68 8.315 2.79 ;
        RECT 6.955 2.2 7.075 2.79 ;
        RECT 4.375 2.29 4.615 2.79 ;
        RECT 3.475 2.05 3.595 2.79 ;
        RECT 2.515 1.73 2.635 2.79 ;
        RECT 1.785 1.34 1.905 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.87 1.675 8.735 1.675 8.735 1.8 8.615 1.8 8.615 1.555 8.75 1.555 8.75 0.9 8.735 0.9 8.735 0.66 8.135 0.66 8.135 0.54 7.515 0.54 7.515 1.46 7.395 1.46 7.395 0.56 5.675 0.56 5.675 1.46 5.555 1.46 5.555 0.56 5.195 0.56 5.195 0.52 5.075 0.52 5.075 0.4 5.315 0.4 5.315 0.44 6.245 0.44 6.245 0.4 6.485 0.4 6.485 0.44 7.395 0.44 7.395 0.42 7.755 0.42 7.755 0.4 7.995 0.4 7.995 0.42 8.255 0.42 8.255 0.54 8.855 0.54 8.855 0.78 8.87 0.78 ;
      POLYGON 7.755 1.7 7.675 1.7 7.675 1.94 6.835 1.94 6.835 2.22 4.735 2.22 4.735 2.17 4.055 2.17 4.055 2.05 4.855 2.05 4.855 2.1 6.715 2.1 6.715 1.82 7.555 1.82 7.555 1.58 7.635 1.58 7.635 0.66 7.755 0.66 ;
      POLYGON 7.195 1.46 7.075 1.46 7.075 1.18 6.245 1.18 6.245 1.62 6.355 1.62 6.355 1.74 6.115 1.74 6.115 1.62 6.125 1.62 6.125 1.26 6.035 1.26 6.035 1.02 6.125 1.02 6.125 0.72 6.365 0.72 6.365 0.84 6.245 0.84 6.245 1.06 7.195 1.06 ;
      POLYGON 6.915 1.42 6.795 1.42 6.795 1.7 6.595 1.7 6.595 1.98 5.785 1.98 5.785 1.96 5.065 1.96 5.065 1.6 4.8 1.6 4.8 1.57 4.135 1.57 4.135 1.69 3.895 1.69 3.895 1.57 4.015 1.57 4.015 1.45 4.275 1.45 4.275 0.66 4.395 0.66 4.395 1.45 4.92 1.45 4.92 1.48 5.185 1.48 5.185 1.84 5.785 1.84 5.785 1.58 5.795 1.58 5.795 0.68 5.915 0.68 5.915 1.7 5.905 1.7 5.905 1.86 6.475 1.86 6.475 1.58 6.675 1.58 6.675 1.3 6.915 1.3 ;
      POLYGON 5.545 1.72 5.305 1.72 5.305 1.16 4.515 1.16 4.515 0.54 4.155 0.54 4.155 0.72 4.035 0.72 4.035 1.08 2.385 1.08 2.385 1.22 2.265 1.22 2.265 0.96 3.915 0.96 3.915 0.6 4.035 0.6 4.035 0.42 4.635 0.42 4.635 1.04 5.305 1.04 5.305 0.86 5.195 0.86 5.195 0.74 5.435 0.74 5.435 0.86 5.425 0.86 5.425 1.6 5.545 1.6 ;
      POLYGON 4.955 0.92 4.835 0.92 4.835 0.6 4.755 0.6 4.755 0.36 4.875 0.36 4.875 0.48 4.955 0.48 ;
      POLYGON 4.945 1.84 4.825 1.84 4.825 1.93 2.995 1.93 2.995 1.63 3.115 1.63 3.115 1.81 4.705 1.81 4.705 1.72 4.945 1.72 ;
      POLYGON 3.915 0.48 3.795 0.48 3.795 0.72 2.775 0.72 2.775 0.84 2.535 0.84 2.535 0.72 2.655 0.72 2.655 0.6 3.675 0.6 3.675 0.36 3.915 0.36 ;
      POLYGON 2.895 1.37 2.625 1.37 2.625 1.46 2.325 1.46 2.325 1.58 2.205 1.58 2.205 1.46 2.025 1.46 2.025 1.2 1.605 1.2 1.605 1.08 2.025 1.08 2.025 0.72 2.385 0.72 2.385 0.84 2.145 0.84 2.145 1.34 2.505 1.34 2.505 1.25 2.895 1.25 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFSX1

MACRO FILL2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL2 0 0 ;
  SIZE 0.58 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.58 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.58 0.18 ;
    END
  END VSS
END FILL2

MACRO DFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRXL 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.945 1.485 2.065 1.75 ;
        RECT 1.81 1.445 1.96 1.725 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.755 2.13 7.635 2.25 ;
        RECT 6.755 1.73 6.875 2.25 ;
        RECT 6.155 1.73 6.875 1.85 ;
        RECT 5.185 1.84 6.275 1.9 ;
        RECT 5.695 1.78 6.875 1.85 ;
        RECT 5.185 1.84 5.815 1.96 ;
        RECT 3.915 1.74 5.305 1.86 ;
        RECT 3.215 1.81 4.035 1.93 ;
        RECT 3.215 1.25 3.455 1.37 ;
        RECT 3.215 1.25 3.335 1.93 ;
        RECT 2.915 1.52 3.335 1.67 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.375 0.87 9.515 1.22 ;
        RECT 9.33 0.81 9.5 1.16 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.2 10.715 1.43 ;
        RECT 10.465 1.2 10.585 1.61 ;
    END
  END CKN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 1.585 1.485 2.09 ;
        RECT 1.365 0.68 1.485 0.96 ;
        RECT 1.23 1.465 1.445 1.725 ;
        RECT 1.325 0.84 1.445 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.765 -0.18 10.885 0.4 ;
        RECT 9.355 -0.18 9.475 0.38 ;
        RECT 8.035 -0.18 8.275 0.33 ;
        RECT 3.075 -0.18 3.315 0.32 ;
        RECT 1.785 -0.18 1.905 0.92 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.705 1.67 10.825 2.79 ;
        RECT 9.315 1.9 9.435 2.79 ;
        RECT 7.775 2.13 7.895 2.79 ;
        RECT 6.175 2.29 6.415 2.79 ;
        RECT 4.415 2.22 4.655 2.79 ;
        RECT 3.075 2.29 3.315 2.79 ;
        RECT 1.785 1.97 1.905 2.79 ;
        RECT 0.555 1.46 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.465 1.85 10.215 1.85 10.215 0.96 10.285 0.96 10.285 0.6 9.715 0.6 9.715 0.62 9.105 0.62 9.105 0.57 7.595 0.57 7.595 0.48 7.475 0.48 7.475 0.36 7.715 0.36 7.715 0.45 8.575 0.45 8.575 0.38 8.815 0.38 8.815 0.45 9.225 0.45 9.225 0.5 9.595 0.5 9.595 0.38 9.915 0.38 9.915 0.48 10.405 0.48 10.405 1.08 10.335 1.08 10.335 1.73 10.465 1.73 ;
      POLYGON 10.075 0.84 9.955 0.84 9.955 1.78 9.875 1.78 9.875 2.02 9.755 2.02 9.755 1.78 9.095 1.78 9.095 2.2 8.375 2.2 8.375 2.01 6.995 2.01 6.995 1.61 6.675 1.61 6.675 1.35 6.245 1.35 6.245 1.23 6.795 1.23 6.795 1.49 7.115 1.49 7.115 1.89 8.495 1.89 8.495 2.08 8.975 2.08 8.975 1.53 8.515 1.53 8.515 1.29 8.635 1.29 8.635 1.41 8.975 1.41 8.975 1.28 9.235 1.28 9.235 1.4 9.095 1.4 9.095 1.66 9.835 1.66 9.835 0.72 10.075 0.72 ;
      POLYGON 8.975 0.84 8.855 0.84 8.855 1.13 8.395 1.13 8.395 1.65 8.735 1.65 8.735 1.84 8.855 1.84 8.855 1.96 8.615 1.96 8.615 1.77 8.275 1.77 8.275 1.13 7.155 1.13 7.155 1.01 8.735 1.01 8.735 0.72 8.975 0.72 ;
      POLYGON 8.155 1.53 7.915 1.53 7.915 1.37 7.355 1.37 7.355 1.65 7.475 1.65 7.475 1.77 7.235 1.77 7.235 1.37 6.915 1.37 6.915 1.11 6.125 1.11 6.125 1.58 6.035 1.58 6.035 1.66 5.785 1.66 5.785 1.54 5.915 1.54 5.915 1.46 6.005 1.46 6.005 0.86 5.885 0.86 5.885 0.62 6.005 0.62 6.005 0.74 6.125 0.74 6.125 0.99 6.915 0.99 6.915 0.75 6.995 0.75 6.995 0.63 7.115 0.63 7.115 0.87 7.035 0.87 7.035 1.25 8.035 1.25 8.035 1.41 8.155 1.41 ;
      POLYGON 7.595 0.81 7.355 0.81 7.355 0.72 7.235 0.72 7.235 0.51 6.695 0.51 6.695 0.87 6.575 0.87 6.575 0.39 7.355 0.39 7.355 0.6 7.475 0.6 7.475 0.69 7.595 0.69 ;
      POLYGON 6.635 2.09 6.515 2.09 6.515 2.14 6.055 2.14 6.055 2.2 4.875 2.2 4.875 2.1 4.275 2.1 4.275 2.22 4.155 2.22 4.155 2.17 2.205 2.17 2.205 1.85 2.265 1.85 2.265 0.68 2.385 0.68 2.385 2.05 4.155 2.05 4.155 1.98 4.995 1.98 4.995 2.08 5.935 2.08 5.935 2.02 6.395 2.02 6.395 1.97 6.635 1.97 ;
      POLYGON 5.885 1.34 5.645 1.34 5.645 0.48 5.205 0.48 5.205 0.36 5.765 0.36 5.765 1.22 5.885 1.22 ;
      POLYGON 5.545 1.72 5.425 1.72 5.425 1.58 5.405 1.58 5.405 1.38 3.575 1.38 3.575 1.13 3.095 1.13 3.095 1.18 2.855 1.18 2.855 1.06 2.975 1.06 2.975 1.01 3.695 1.01 3.695 1.26 5.405 1.26 5.405 0.62 5.525 0.62 5.525 1.46 5.545 1.46 ;
      POLYGON 5.185 1.62 3.795 1.62 3.795 1.69 3.555 1.69 3.555 1.57 3.675 1.57 3.675 1.5 5.185 1.5 ;
      POLYGON 5.105 0.86 4.955 0.86 4.955 1.14 4.355 1.14 4.355 0.9 4.175 0.9 4.175 0.66 4.295 0.66 4.295 0.78 4.475 0.78 4.475 1.02 4.835 1.02 4.835 0.74 4.985 0.74 4.985 0.62 5.105 0.62 ;
      POLYGON 4.715 0.9 4.595 0.9 4.595 0.54 4.055 0.54 4.055 0.76 3.795 0.76 3.795 0.84 3.555 0.84 3.555 0.72 3.675 0.72 3.675 0.64 3.935 0.64 3.935 0.42 4.715 0.42 ;
      POLYGON 3.815 0.52 3.555 0.52 3.555 0.56 2.775 0.56 2.775 0.9 2.735 0.9 2.735 1.3 2.775 1.3 2.775 1.75 2.655 1.75 2.655 1.42 2.615 1.42 2.615 0.78 2.655 0.78 2.655 0.56 2.145 0.56 2.145 1.2 1.565 1.2 1.565 1.08 2.025 1.08 2.025 0.44 3.435 0.44 3.435 0.4 3.815 0.4 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFNSRXL

MACRO OAI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X4 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.305 1.26 5.085 1.38 ;
        RECT 4.365 1.23 4.625 1.38 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.065 1.2 6.705 1.32 ;
        RECT 6.585 1.08 6.705 1.32 ;
        RECT 6.45 1.175 6.6 1.435 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.195 1.04 3.435 1.16 ;
        RECT 0.68 0.99 3.315 1.11 ;
        RECT 1.835 0.99 2.075 1.16 ;
        RECT 0.65 1.02 0.8 1.435 ;
        RECT 0.435 1.02 0.8 1.14 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.28 2.715 1.4 ;
        RECT 2.335 1.23 2.595 1.4 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.825 0.81 6.965 0.93 ;
        RECT 6.845 0.64 6.965 0.93 ;
        RECT 6.605 1.555 6.725 2.21 ;
        RECT 1.415 1.555 6.725 1.675 ;
        RECT 5.825 0.76 6.125 0.93 ;
        RECT 6.005 0.64 6.125 0.93 ;
        RECT 4.065 0.99 5.945 1.11 ;
        RECT 5.825 0.76 5.945 1.11 ;
        RECT 5.765 1.555 5.885 2.21 ;
        RECT 4.925 1.555 5.045 2.21 ;
        RECT 4.065 1.52 4.335 1.675 ;
        RECT 4.085 1.52 4.205 2.21 ;
        RECT 4.065 0.99 4.185 1.675 ;
        RECT 2.695 1.555 2.815 2.21 ;
        RECT 1.415 1.555 1.535 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 3.455 0.51 3.695 0.63 ;
        RECT 3.455 -0.18 3.575 0.63 ;
        RECT 2.615 0.51 2.855 0.63 ;
        RECT 2.615 -0.18 2.735 0.63 ;
        RECT 1.775 0.51 2.015 0.63 ;
        RECT 1.775 -0.18 1.895 0.63 ;
        RECT 0.935 0.51 1.175 0.63 ;
        RECT 0.935 -0.18 1.055 0.63 ;
        RECT 0.155 -0.18 0.275 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 7.025 1.56 7.145 2.79 ;
        RECT 6.185 1.795 6.305 2.79 ;
        RECT 5.345 1.795 5.465 2.79 ;
        RECT 4.445 1.795 4.685 2.15 ;
        RECT 4.445 1.795 4.565 2.79 ;
        RECT 3.665 1.795 3.785 2.79 ;
        RECT 2.055 1.795 2.175 2.79 ;
        RECT 0.355 1.56 0.475 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.385 0.69 7.265 0.69 7.265 0.52 6.545 0.52 6.545 0.69 6.425 0.69 6.425 0.52 5.705 0.52 5.705 0.69 5.585 0.69 5.585 0.52 4.925 0.52 4.925 0.63 4.685 0.63 4.685 0.52 4.085 0.52 4.085 0.63 3.845 0.63 3.845 0.51 3.965 0.51 3.965 0.4 7.385 0.4 ;
      POLYGON 5.345 0.82 5.225 0.82 5.225 0.87 0.575 0.87 0.575 0.63 0.695 0.63 0.695 0.75 1.415 0.75 1.415 0.63 1.535 0.63 1.535 0.75 2.255 0.75 2.255 0.63 2.375 0.63 2.375 0.75 3.095 0.75 3.095 0.63 3.215 0.63 3.215 0.75 4.265 0.75 4.265 0.7 4.505 0.7 4.505 0.75 5.105 0.75 5.105 0.7 5.345 0.7 ;
  END
END OAI211X4

MACRO TLATNCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX8 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.465 0.565 1.67 ;
        RECT 0.445 1.26 0.565 1.67 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.515 1.145 1.72 ;
        RECT 0.915 1.36 1.035 1.72 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.155 1.1 8.275 2.08 ;
        RECT 8.135 0.645 8.255 1.22 ;
        RECT 5.61 1.1 8.275 1.22 ;
        RECT 6.515 0.765 8.255 0.885 ;
        RECT 7.235 0.715 7.475 0.885 ;
        RECT 7.315 1.1 7.435 2.08 ;
        RECT 6.395 0.715 6.635 0.835 ;
        RECT 6.475 1.1 6.595 2.085 ;
        RECT 5.635 1.1 5.755 2.085 ;
        RECT 5.555 0.885 5.73 1.1 ;
        RECT 5.555 0.655 5.675 1.1 ;
        RECT 5.61 1.1 5.755 1.34 ;
        RECT 5.58 1.1 8.275 1.145 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.715 -0.18 7.835 0.645 ;
        RECT 6.875 -0.18 6.995 0.645 ;
        RECT 5.975 -0.18 6.095 0.64 ;
        RECT 5.135 -0.18 5.255 0.64 ;
        RECT 3.735 0.45 3.975 0.57 ;
        RECT 3.855 -0.18 3.975 0.57 ;
        RECT 2.275 -0.18 2.395 0.38 ;
        RECT 0.555 -0.18 0.675 0.9 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.735 1.34 7.855 2.79 ;
        RECT 6.895 1.34 7.015 2.79 ;
        RECT 6.055 1.34 6.175 2.79 ;
        RECT 5.215 1.77 5.335 2.79 ;
        RECT 4.375 1.77 4.495 2.79 ;
        RECT 3.475 2.23 3.595 2.79 ;
        RECT 2.075 2.26 2.315 2.79 ;
        RECT 0.755 1.84 0.875 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.435 1.215 5.335 1.215 5.335 1.65 4.915 1.65 4.915 2.08 4.795 2.08 4.795 1.65 4.075 1.65 4.075 2.08 3.955 2.08 3.955 1.53 5.215 1.53 5.215 0.97 4.575 0.97 4.575 0.81 4.495 0.81 4.495 0.57 4.615 0.57 4.615 0.69 4.695 0.69 4.695 0.85 5.435 0.85 ;
      POLYGON 5.095 1.41 3.875 1.41 3.875 1.05 3.255 1.05 3.255 1.43 3.125 1.43 3.125 1.87 3.005 1.87 3.005 1.43 2.075 1.43 2.075 1.31 3.135 1.31 3.135 0.65 3.375 0.65 3.375 0.77 3.255 0.77 3.255 0.93 3.995 0.93 3.995 1.29 4.975 1.29 4.975 1.09 5.095 1.09 ;
      POLYGON 4.455 1.17 4.335 1.17 4.335 1.05 4.255 1.05 4.255 0.81 3.495 0.81 3.495 0.53 3.015 0.53 3.015 0.74 2.875 0.74 2.875 1.18 1.955 1.18 1.955 1.74 2.675 1.74 2.675 1.78 2.795 1.78 2.795 1.9 2.555 1.9 2.555 1.86 1.835 1.86 1.835 1.18 1.755 1.18 1.755 1.06 2.755 1.06 2.755 0.62 2.895 0.62 2.895 0.41 3.615 0.41 3.615 0.69 4.375 0.69 4.375 0.93 4.455 0.93 ;
      POLYGON 3.615 1.29 3.495 1.29 3.495 2.11 3.145 2.11 3.145 2.14 2.23 2.14 2.23 2.1 1.435 2.1 1.435 1.86 1.275 1.86 1.275 0.66 1.395 0.66 1.395 1.74 1.555 1.74 1.555 1.98 2.35 1.98 2.35 2.02 3.025 2.02 3.025 1.99 3.375 1.99 3.375 1.17 3.615 1.17 ;
      POLYGON 2.775 0.5 2.635 0.5 2.635 0.62 2.035 0.62 2.035 0.54 1.635 0.54 1.635 1.38 1.715 1.38 1.715 1.62 1.515 1.62 1.515 0.54 1.155 0.54 1.155 1.24 1.035 1.24 1.035 1.14 0.185 1.14 0.185 1.79 0.455 1.79 0.455 2.03 0.335 2.03 0.335 1.91 0.065 1.91 0.065 0.9 0.135 0.9 0.135 0.66 0.255 0.66 0.255 1.02 1.035 1.02 1.035 0.42 2.155 0.42 2.155 0.5 2.515 0.5 2.515 0.38 2.775 0.38 ;
  END
END TLATNCAX8

MACRO BUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX12 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.45 1.3 4.775 1.42 ;
        RECT 4.42 1.465 4.57 1.725 ;
        RECT 4.45 1.3 4.57 1.725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.915 1.32 4.035 2.21 ;
        RECT 0.515 0.82 4.035 0.94 ;
        RECT 3.915 0.4 4.035 0.94 ;
        RECT 0.515 1.32 4.035 1.44 ;
        RECT 3.075 1.32 3.195 2.21 ;
        RECT 3.075 0.4 3.195 0.94 ;
        RECT 2.235 1.32 2.355 2.21 ;
        RECT 2.235 0.4 2.355 0.94 ;
        RECT 1.395 1.32 1.515 2.21 ;
        RECT 1.395 0.4 1.515 0.94 ;
        RECT 0.555 1.32 0.8 1.725 ;
        RECT 0.555 1.32 0.675 2.21 ;
        RECT 0.555 0.4 0.675 0.94 ;
        RECT 0.515 0.8 0.635 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.175 -0.18 5.295 0.725 ;
        RECT 4.335 -0.18 4.455 0.915 ;
        RECT 3.495 -0.18 3.615 0.7 ;
        RECT 2.655 -0.18 2.775 0.7 ;
        RECT 1.815 -0.18 1.935 0.7 ;
        RECT 0.975 -0.18 1.095 0.7 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.175 1.56 5.295 2.79 ;
        RECT 4.335 1.845 4.455 2.79 ;
        RECT 3.495 1.56 3.615 2.79 ;
        RECT 2.655 1.56 2.775 2.79 ;
        RECT 1.815 1.56 1.935 2.79 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.43 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.715 0.965 5.015 0.965 5.015 1.32 5.715 1.32 5.715 2.21 5.595 2.21 5.595 1.44 5.015 1.44 5.015 1.66 4.875 1.66 4.875 2.21 4.755 2.21 4.755 1.54 4.895 1.54 4.895 1.18 3.935 1.18 3.935 1.195 3.695 1.195 3.695 1.18 3.095 1.18 3.095 1.195 2.855 1.195 2.855 1.18 2.675 1.18 2.675 1.195 2.435 1.195 2.435 1.18 1.835 1.18 1.835 1.195 1.595 1.195 1.595 1.18 0.995 1.18 0.995 1.2 0.755 1.2 0.755 1.08 0.875 1.08 0.875 1.06 4.755 1.06 4.755 0.675 4.875 0.675 4.875 0.845 5.595 0.845 5.595 0.675 5.715 0.675 ;
  END
END BUFX12

MACRO AOI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X4 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.715 0.99 6.675 1.11 ;
        RECT 3.785 0.94 4.045 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.99 3.355 1.18 ;
        RECT 3.235 0.94 3.355 1.18 ;
        RECT 2.97 0.99 3.12 1.435 ;
        RECT 0.435 0.99 3.355 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.23 2.775 1.35 ;
        RECT 1.465 1.23 1.725 1.38 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.355 1.26 5.875 1.38 ;
        RECT 5.525 1.23 5.785 1.38 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 1.5 6.555 2.01 ;
        RECT 3.915 1.5 6.555 1.62 ;
        RECT 5.595 1.5 5.715 2.01 ;
        RECT 5.475 0.65 5.715 0.77 ;
        RECT 1.535 0.7 5.595 0.82 ;
        RECT 4.755 1.5 4.875 2.01 ;
        RECT 4.195 0.65 4.435 0.82 ;
        RECT 3.915 1.315 4.035 2.01 ;
        RECT 3.475 1.315 4.035 1.435 ;
        RECT 3.475 1.23 3.755 1.435 ;
        RECT 3.475 0.7 3.595 1.435 ;
        RECT 2.695 0.65 2.935 0.82 ;
        RECT 1.415 0.65 1.655 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.175 -0.18 6.295 0.64 ;
        RECT 4.835 0.46 5.075 0.58 ;
        RECT 4.835 -0.18 4.955 0.58 ;
        RECT 3.435 0.46 3.675 0.58 ;
        RECT 3.435 -0.18 3.555 0.58 ;
        RECT 2.055 0.46 2.295 0.58 ;
        RECT 2.055 -0.18 2.175 0.58 ;
        RECT 0.835 -0.18 0.955 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 3.075 1.795 3.195 2.79 ;
        RECT 2.235 1.795 2.355 2.79 ;
        RECT 1.395 1.795 1.515 2.79 ;
        RECT 0.555 1.795 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.975 2.25 3.495 2.25 3.495 1.675 2.775 1.675 2.775 2.21 2.655 2.21 2.655 1.675 1.935 1.675 1.935 2.21 1.815 2.21 1.815 1.675 1.095 1.675 1.095 2.21 0.975 2.21 0.975 1.675 0.255 1.675 0.255 2.21 0.135 2.21 0.135 1.555 3.615 1.555 3.615 2.13 4.335 2.13 4.335 1.74 4.455 1.74 4.455 2.13 5.175 2.13 5.175 1.74 5.295 1.74 5.295 2.13 6.015 2.13 6.015 1.74 6.135 1.74 6.135 2.13 6.855 2.13 6.855 1.56 6.975 1.56 ;
  END
END AOI22X4

MACRO OAI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X2 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.075 0.66 8.375 0.78 ;
        RECT 8.255 0.54 8.375 0.78 ;
        RECT 7.355 0.855 8.195 0.975 ;
        RECT 8.075 0.66 8.195 0.975 ;
        RECT 1.455 1.845 7.995 1.965 ;
        RECT 7.875 0.855 7.995 1.965 ;
        RECT 7.355 0.6 7.595 0.72 ;
        RECT 4.82 0.79 7.475 0.91 ;
        RECT 7.355 0.6 7.475 0.975 ;
        RECT 6.455 0.6 6.695 0.91 ;
        RECT 5.615 0.6 5.855 0.91 ;
        RECT 4.655 0.65 5.015 0.8 ;
        RECT 4.775 0.6 5.015 0.8 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.97 2.815 1.09 ;
        RECT 2.335 0.94 2.595 1.09 ;
    END
  END A0
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.74 1.03 7.175 1.15 ;
        RECT 4.74 1.03 4.955 1.295 ;
        RECT 4.71 1.175 4.86 1.435 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.23 3.775 1.35 ;
        RECT 3.495 1.23 3.755 1.38 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.135 1.27 7.495 1.39 ;
        RECT 5.135 1.27 5.255 1.535 ;
        RECT 5 1.465 5.215 1.655 ;
        RECT 5 1.465 5.15 1.725 ;
        RECT 5.03 1.415 5.255 1.535 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 1.52 4.335 1.67 ;
        RECT 1.295 1.5 4.315 1.61 ;
        RECT 4.075 1.49 4.315 1.67 ;
        RECT 1.945 1.52 4.335 1.62 ;
        RECT 1.295 1.49 2.065 1.61 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.635 1.44 7.755 1.68 ;
        RECT 5.475 1.51 7.755 1.63 ;
        RECT 5.525 1.51 5.785 1.67 ;
    END
  END B0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 3.855 0.46 4.095 0.58 ;
        RECT 3.855 -0.18 3.975 0.58 ;
        RECT 2.895 0.46 3.135 0.58 ;
        RECT 2.895 -0.18 3.015 0.58 ;
        RECT 1.935 0.46 2.175 0.58 ;
        RECT 1.935 -0.18 2.055 0.58 ;
        RECT 0.975 0.46 1.215 0.58 ;
        RECT 0.975 -0.18 1.095 0.58 ;
        RECT 0.135 -0.18 0.255 0.725 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.795 2.085 8.035 2.205 ;
        RECT 7.795 2.085 7.915 2.79 ;
        RECT 5.655 2.085 5.895 2.205 ;
        RECT 5.655 2.085 5.775 2.79 ;
        RECT 2.475 2.085 2.715 2.205 ;
        RECT 2.475 2.085 2.595 2.79 ;
        RECT 0.335 1.97 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.955 0.735 7.835 0.735 7.835 0.48 7.115 0.48 7.115 0.67 6.875 0.67 6.875 0.48 6.275 0.48 6.275 0.67 6.035 0.67 6.035 0.48 5.435 0.48 5.435 0.67 5.195 0.67 5.195 0.48 4.535 0.48 4.535 0.82 0.555 0.82 0.555 0.535 0.675 0.535 0.675 0.7 1.515 0.7 1.515 0.535 1.635 0.535 1.635 0.7 2.475 0.7 2.475 0.535 2.595 0.535 2.595 0.7 3.435 0.7 3.435 0.535 3.555 0.535 3.555 0.7 4.415 0.7 4.415 0.36 7.955 0.36 ;
  END
END OAI33X2

MACRO EDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX2 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.23 0.855 1.4 ;
        RECT 0.47 1.23 0.855 1.385 ;
        RECT 0.47 1.11 0.59 1.385 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.82 1.13 8.06 1.335 ;
        RECT 7.9 1.08 8.05 1.475 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.19 0.84 8.34 1.145 ;
        RECT 7.16 0.84 8.34 0.96 ;
        RECT 7.32 0.36 7.44 0.96 ;
        RECT 6.68 0.36 7.44 0.48 ;
        RECT 7.16 0.84 7.28 1.17 ;
        RECT 6.68 0.36 6.8 1.27 ;
        RECT 6.58 1.15 6.7 1.39 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.42 1.53 5.66 1.65 ;
        RECT 5.42 0.67 5.66 0.79 ;
        RECT 5.42 0.67 5.54 1.65 ;
        RECT 5.29 1.175 5.54 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.66 -0.18 7.78 0.66 ;
        RECT 6.02 -0.18 6.14 0.66 ;
        RECT 4.94 -0.18 5.06 0.68 ;
        RECT 2.96 0.49 3.2 0.61 ;
        RECT 2.96 -0.18 3.08 0.61 ;
        RECT 0.59 0.57 0.83 0.69 ;
        RECT 0.59 -0.18 0.71 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 8.02 1.835 8.14 2.79 ;
        RECT 5.9 2.01 6.14 2.13 ;
        RECT 5.9 2.01 6.02 2.79 ;
        RECT 4.94 2.01 5.18 2.13 ;
        RECT 4.94 2.01 5.06 2.79 ;
        RECT 3.02 1.72 3.14 2.79 ;
        RECT 2.9 1.72 3.14 1.93 ;
        RECT 0.65 1.57 0.77 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.58 1.835 8.56 1.835 8.56 2 8.44 2 8.44 1.715 7.52 1.715 7.52 1.15 7.64 1.15 7.64 1.595 8.46 1.595 8.46 0.72 8.38 0.72 8.38 0.48 8.5 0.48 8.5 0.6 8.58 0.6 ;
      POLYGON 7.2 0.72 7.04 0.72 7.04 2.12 6.92 2.12 6.92 1.89 4.705 1.89 4.705 2.23 3.26 2.23 3.26 1.6 2.78 1.6 2.78 2.23 1.66 2.23 1.66 1.59 1.5 1.59 1.5 0.72 1.4 0.72 1.4 0.6 1.64 0.6 1.64 0.72 1.62 0.72 1.62 1.47 1.78 1.47 1.78 2.11 2.66 2.11 2.66 1.48 3.38 1.48 3.38 2.11 4.585 2.11 4.585 1.77 6.92 1.77 6.92 0.6 7.2 0.6 ;
      POLYGON 6.62 1.65 6.34 1.65 6.34 1.41 5.74 1.41 5.74 1.15 5.86 1.15 5.86 1.29 6.34 1.29 6.34 0.73 6.44 0.73 6.44 0.61 6.56 0.61 6.56 0.85 6.46 0.85 6.46 1.53 6.62 1.53 ;
      POLYGON 6.22 1.17 6.1 1.17 6.1 0.9 5.78 0.9 5.78 0.55 5.3 0.55 5.3 0.92 4.8 0.92 4.8 1.63 4.32 1.63 4.32 1.99 4.2 1.99 4.2 1.47 4.32 1.47 4.32 1.51 4.68 1.51 4.68 0.92 4.16 0.92 4.16 0.54 4.28 0.54 4.28 0.8 5.18 0.8 5.18 0.43 5.9 0.43 5.9 0.78 6.22 0.78 ;
      POLYGON 4.56 1.39 4.44 1.39 4.44 1.16 3.92 1.16 3.92 1.04 3.8 1.04 3.8 0.92 3.92 0.92 3.92 0.48 3.44 0.48 3.44 0.85 2.625 0.85 2.625 0.48 2.48 0.48 2.48 1.12 2.36 1.12 2.36 0.48 1.88 0.48 1.88 1.21 1.98 1.21 1.98 1.33 1.74 1.33 1.74 1.21 1.76 1.21 1.76 0.48 1.19 0.48 1.19 0.63 1.23 0.63 1.23 1.57 1.19 1.57 1.19 1.69 1.07 1.69 1.07 1.45 1.11 1.45 1.11 0.75 1.07 0.75 1.07 0.36 2.745 0.36 2.745 0.73 3.32 0.73 3.32 0.36 4.04 0.36 4.04 1.04 4.56 1.04 ;
      POLYGON 3.8 0.72 3.68 0.72 3.68 1.33 3.62 1.33 3.62 1.99 3.5 1.99 3.5 1.33 2.84 1.33 2.84 1.21 3.56 1.21 3.56 0.6 3.8 0.6 ;
      POLYGON 3.44 1.09 2.72 1.09 2.72 1.36 2.24 1.36 2.24 1.99 2.12 1.99 2.12 0.72 2 0.72 2 0.6 2.24 0.6 2.24 1.24 2.6 1.24 2.6 0.97 3.44 0.97 ;
      POLYGON 0.99 1.01 0.75 1.01 0.75 0.99 0.35 0.99 0.35 1.69 0.23 1.69 0.23 0.51 0.35 0.51 0.35 0.87 0.99 0.87 ;
  END
END EDFFHQX2

MACRO AND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.065 0.51 1.46 ;
        RECT 0.24 1.09 0.51 1.295 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.93 0.82 1.355 ;
        RECT 0.65 1.055 0.8 1.46 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 0.93 1.16 1.28 ;
        RECT 0.94 1.11 1.09 1.46 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.575 1.02 1.695 1.46 ;
        RECT 1.52 1.02 1.695 1.44 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.355 1.34 2.475 1.99 ;
        RECT 2.045 1.23 2.435 1.38 ;
        RECT 2.315 0.73 2.435 1.46 ;
        RECT 2.215 0.61 2.335 0.85 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.795 -0.18 1.915 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.935 1.5 2.055 2.79 ;
        RECT 1.035 2.14 1.155 2.79 ;
        RECT 0.135 1.62 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.195 1.11 1.955 1.11 1.955 0.9 1.4 0.9 1.4 1.58 1.635 1.58 1.635 1.82 1.515 1.82 1.515 1.7 0.495 1.7 0.495 1.58 1.28 1.58 1.28 0.81 0.28 0.81 0.28 0.79 0.16 0.79 0.16 0.67 0.4 0.67 0.4 0.69 1.4 0.69 1.4 0.78 2.075 0.78 2.075 0.99 2.195 0.99 ;
  END
END AND4X1

MACRO CLKMX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X8 0 0 ;
  SIZE 5.8 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.12 1.505 1.24 ;
        RECT 0.645 1.5 1.385 1.62 ;
        RECT 1.265 1.12 1.385 1.62 ;
        RECT 0.645 1.175 0.765 1.62 ;
        RECT 0.36 1.175 0.765 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.11 1.145 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.08 2.54 1.46 ;
        RECT 2.28 1.08 2.54 1.275 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.725 0.765 5.465 0.885 ;
        RECT 5.345 0.645 5.465 0.885 ;
        RECT 5.34 0.765 5.46 2.205 ;
        RECT 2.97 1.225 5.46 1.345 ;
        RECT 4.445 0.715 4.685 0.885 ;
        RECT 4.5 1.225 4.62 2.205 ;
        RECT 3.605 0.715 3.845 0.835 ;
        RECT 3.66 1.225 3.78 2.21 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 2.82 1.345 3.09 1.465 ;
        RECT 2.97 0.6 3.09 1.465 ;
        RECT 2.765 0.6 3.09 0.72 ;
        RECT 2.82 1.345 2.94 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.8 0.18 ;
        RECT 4.925 -0.18 5.045 0.645 ;
        RECT 4.085 -0.18 4.205 0.645 ;
        RECT 3.245 -0.18 3.365 0.645 ;
        RECT 2.345 0.46 2.585 0.58 ;
        RECT 2.345 -0.18 2.465 0.58 ;
        RECT 0.825 -0.18 0.945 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.8 2.79 ;
        RECT 4.92 1.465 5.04 2.79 ;
        RECT 4.08 1.465 4.2 2.79 ;
        RECT 3.24 1.465 3.36 2.79 ;
        RECT 2.4 1.58 2.52 2.79 ;
        RECT 0.96 1.74 1.2 2.14 ;
        RECT 0.96 1.74 1.08 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.8 1.215 2.68 1.215 2.68 0.96 2.16 0.96 2.16 1.78 1.78 1.78 1.78 2.2 1.66 2.2 1.66 1.66 2.04 1.66 2.04 0.96 1.985 0.96 1.985 0.75 1.765 0.75 1.765 0.5 1.885 0.5 1.885 0.63 2.105 0.63 2.105 0.84 2.8 0.84 ;
      POLYGON 1.92 1.54 1.625 1.54 1.625 0.99 0.24 0.99 0.24 1.555 0.525 1.555 0.525 1.92 0.405 1.92 0.405 1.675 0.12 1.675 0.12 0.75 0.345 0.75 0.345 0.5 0.465 0.5 0.465 0.87 1.745 0.87 1.745 0.88 1.865 0.88 1.865 1 1.745 1 1.745 1.42 1.92 1.42 ;
  END
END CLKMX2X8

MACRO MXI2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 1.335 1.74 1.455 ;
        RECT 1.62 1.135 1.74 1.455 ;
        RECT 0.99 1.335 1.18 1.575 ;
        RECT 0.39 1.555 1.11 1.675 ;
        RECT 0.39 1.175 0.51 1.675 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 1.175 0.87 1.435 ;
        RECT 0.65 1.135 0.87 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.135 2.32 1.44 ;
        RECT 2.1 1.135 2.295 1.46 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.6 1.175 2.83 1.435 ;
        RECT 2.6 0.8 2.72 2.21 ;
        RECT 2.55 0.68 2.67 0.92 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.03 -0.18 3.15 0.38 ;
        RECT 2.07 -0.18 2.19 0.775 ;
        RECT 0.68 -0.18 0.8 0.775 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.02 1.56 3.14 2.79 ;
        RECT 2.18 1.58 2.3 2.79 ;
        RECT 0.58 1.795 0.7 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.69 0.86 3.57 0.86 3.57 1.195 3.63 1.195 3.63 1.8 3.51 1.8 3.51 1.315 2.95 1.315 2.95 1.195 3.45 1.195 3.45 0.74 3.69 0.74 ;
      POLYGON 3.53 0.52 3.41 0.52 3.41 0.62 2.79 0.62 2.79 0.56 2.43 0.56 2.43 1.015 1.98 1.015 1.98 1.695 1.42 1.695 1.42 1.815 1.35 1.815 1.35 1.935 1.23 1.935 1.23 1.695 1.3 1.695 1.3 1.575 1.86 1.575 1.86 1.015 1.595 1.015 1.595 0.775 1.43 0.775 1.43 0.535 1.55 0.535 1.55 0.655 1.715 0.655 1.715 0.895 2.31 0.895 2.31 0.44 2.91 0.44 2.91 0.5 3.29 0.5 3.29 0.4 3.53 0.4 ;
      POLYGON 1.29 1.135 1.17 1.135 1.17 1.015 0.24 1.015 0.24 1.795 0.28 1.795 0.28 2.035 0.16 2.035 0.16 1.915 0.12 1.915 0.12 0.775 0.26 0.775 0.26 0.535 0.38 0.535 0.38 0.895 1.29 0.895 ;
  END
END MXI2X2

MACRO SEDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX1 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.085 0.5 2.205 1.49 ;
        RECT 1.945 0.5 2.205 0.62 ;
        RECT 1.165 0.42 2.065 0.54 ;
        RECT 1.265 0.98 1.385 1.22 ;
        RECT 1.165 0.42 1.285 1.1 ;
        RECT 0.535 0.98 1.385 1.1 ;
        RECT 0.305 1.23 0.655 1.38 ;
        RECT 0.535 0.94 0.655 1.38 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.22 1.145 1.41 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.94 1.055 4.085 1.295 ;
        RECT 3.84 1.175 4.01 1.435 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 0.81 5.73 1.265 ;
        RECT 5.59 0.81 5.71 1.53 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.09 1.085 11.31 1.435 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.71 1.57 3.23 1.69 ;
        RECT 2.71 0.72 2.83 1.69 ;
        RECT 2.665 0.6 2.785 0.84 ;
        RECT 2.68 1.175 2.83 1.435 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.33 1.62 6.57 1.865 ;
        RECT 6.33 0.76 6.45 1.865 ;
        RECT 6.105 0.76 6.45 1.09 ;
        RECT 6.105 0.64 6.225 1.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.03 -0.18 11.15 0.725 ;
        RECT 9.04 0.31 9.28 0.43 ;
        RECT 9.04 -0.18 9.16 0.43 ;
        RECT 7.3 0.45 7.54 0.57 ;
        RECT 7.3 -0.18 7.42 0.57 ;
        RECT 5.625 -0.18 5.745 0.69 ;
        RECT 3.695 -0.18 3.815 0.92 ;
        RECT 2.185 -0.18 2.305 0.38 ;
        RECT 0.725 0.66 0.965 0.78 ;
        RECT 0.845 -0.18 0.965 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 11.09 1.795 11.21 2.79 ;
        RECT 8.92 2.29 9.16 2.79 ;
        RECT 7.26 2.15 7.38 2.79 ;
        RECT 5.85 2.225 6.09 2.79 ;
        RECT 3.86 2.29 4.1 2.79 ;
        RECT 2.57 2.23 2.69 2.79 ;
        RECT 0.725 1.77 0.965 1.89 ;
        RECT 0.725 1.77 0.845 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.69 1.855 11.45 1.855 11.45 1.675 10.97 1.675 10.97 2.23 9.46 2.23 9.46 2.17 8.16 2.17 8.16 2.05 9.7 2.05 9.7 2.11 10.85 2.11 10.85 0.845 11.27 0.845 11.27 0.605 11.45 0.605 11.45 0.485 11.57 0.485 11.57 0.725 11.39 0.725 11.39 0.965 10.97 0.965 10.97 1.555 11.57 1.555 11.57 1.735 11.69 1.735 ;
      POLYGON 10.73 1.99 9.98 1.99 9.98 1.93 8.26 1.93 8.26 1.29 7.92 1.29 7.92 1.41 7.8 1.41 7.8 1.17 8.26 1.17 8.26 1.03 8.54 1.03 8.54 1.15 8.38 1.15 8.38 1.81 9.98 1.81 9.98 1.41 9.94 1.41 9.94 1.17 10.06 1.17 10.06 1.29 10.1 1.29 10.1 1.87 10.61 1.87 10.61 0.485 10.73 0.485 ;
      POLYGON 10.34 1.75 10.22 1.75 10.22 0.48 9.545 0.48 9.545 0.67 8.8 0.67 8.8 0.48 7.78 0.48 7.78 0.81 7.06 0.81 7.06 0.48 5.985 0.48 5.985 1.1 5.97 1.1 5.97 1.865 5.33 1.865 5.33 1.985 5.21 1.985 5.21 1.865 5.1 1.865 5.1 0.88 4.925 0.88 4.925 0.64 5.045 0.64 5.045 0.76 5.22 0.76 5.22 1.745 5.85 1.745 5.85 0.98 5.865 0.98 5.865 0.36 7.18 0.36 7.18 0.69 7.66 0.69 7.66 0.36 8.92 0.36 8.92 0.55 9.425 0.55 9.425 0.36 10.34 0.36 ;
      POLYGON 9.98 0.72 9.82 0.72 9.82 1.57 9.86 1.57 9.86 1.69 9.62 1.69 9.62 1.57 9.7 1.57 9.7 1.37 8.9 1.37 8.9 1.25 9.7 1.25 9.7 0.6 9.98 0.6 ;
      POLYGON 9.42 1.13 9.3 1.13 9.3 1.03 8.78 1.03 8.78 1.69 8.5 1.69 8.5 1.57 8.66 1.57 8.66 0.91 8.44 0.91 8.44 0.6 8.68 0.6 8.68 0.79 8.78 0.79 8.78 0.91 9.3 0.91 9.3 0.89 9.42 0.89 ;
      POLYGON 8.26 0.72 8.02 0.72 8.02 1.05 7.68 1.05 7.68 1.53 8.02 1.53 8.02 1.57 8.14 1.57 8.14 1.69 7.9 1.69 7.9 1.65 7.56 1.65 7.56 1.37 6.98 1.37 6.98 1.25 7.56 1.25 7.56 0.93 7.9 0.93 7.9 0.6 8.26 0.6 ;
      POLYGON 7.44 1.05 6.86 1.05 6.86 1.63 6.9 1.63 6.9 2.105 5.73 2.105 5.73 2.225 4.455 2.225 4.455 2.17 3.54 2.17 3.54 2.05 4.575 2.05 4.575 2.105 5.61 2.105 5.61 1.985 6.09 1.985 6.09 1.22 6.21 1.22 6.21 1.985 6.78 1.985 6.78 1.75 6.74 1.75 6.74 0.72 6.7 0.72 6.7 0.6 6.94 0.6 6.94 0.72 6.86 0.72 6.86 0.93 7.44 0.93 ;
      POLYGON 5.47 1.625 5.35 1.625 5.35 1.505 5.34 1.505 5.34 0.52 4.235 0.52 4.235 0.8 4.325 0.8 4.325 1.45 4.52 1.45 4.52 1.69 4.4 1.69 4.4 1.57 4.205 1.57 4.205 0.92 4.115 0.92 4.115 0.4 4.705 0.4 4.705 0.36 4.945 0.36 4.945 0.4 5.46 0.4 5.46 1.385 5.47 1.385 ;
      POLYGON 4.91 1.945 4.79 1.945 4.79 1.93 1.885 1.93 1.885 1.73 1.845 1.73 1.845 0.86 1.405 0.86 1.405 0.66 1.645 0.66 1.645 0.74 1.965 0.74 1.965 1.61 2.005 1.61 2.005 1.81 4.685 1.81 4.685 0.82 4.445 0.82 4.445 0.7 4.805 0.7 4.805 1.705 4.91 1.705 ;
      POLYGON 3.56 1.69 3.44 1.69 3.44 0.92 3.275 0.92 3.275 0.68 3.01 0.68 3.01 0.48 2.545 0.48 2.545 1.16 2.425 1.16 2.425 0.36 3.13 0.36 3.13 0.56 3.395 0.56 3.395 0.8 3.56 0.8 ;
      POLYGON 1.725 1.65 0.485 1.65 0.485 1.83 0.365 1.83 0.365 1.71 0.065 1.71 0.065 0.99 0.295 0.99 0.295 0.6 0.415 0.6 0.415 1.11 0.185 1.11 0.185 1.53 1.605 1.53 1.605 1.27 1.725 1.27 ;
  END
END SEDFFX1

MACRO SMDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX4 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 1.53 2.235 1.65 ;
        RECT 1.855 0.66 1.975 0.9 ;
        RECT 1.835 0.78 1.955 1.65 ;
        RECT 0.94 1.315 1.955 1.435 ;
        RECT 1.035 1.315 1.275 1.65 ;
        RECT 0.94 1.175 1.155 1.435 ;
        RECT 1.035 0.78 1.155 1.65 ;
        RECT 1.015 0.66 1.135 0.9 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.02 0.51 1.47 ;
        RECT 0.375 0.915 0.495 1.47 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.32 1.06 7.525 1.44 ;
        RECT 7.405 1.05 7.525 1.44 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.06 0.8 9.21 1.2 ;
        RECT 9.04 0.825 9.16 1.24 ;
    END
  END SE
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.38 0.76 9.5 1.24 ;
        RECT 9.35 0.76 9.5 1.215 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.21 10.94 1.345 ;
        RECT 10.455 1.21 10.715 1.38 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.08 0.97 11.2 1.21 ;
        RECT 9.975 0.97 11.2 1.09 ;
        RECT 10.745 0.94 11.005 1.09 ;
        RECT 9.975 0.97 10.095 1.32 ;
        RECT 9.86 1.2 9.98 1.44 ;
    END
  END S0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.92 -0.18 11.04 0.82 ;
        RECT 9.495 -0.18 9.615 0.64 ;
        RECT 7.505 -0.18 7.625 0.81 ;
        RECT 5.275 -0.18 5.515 0.37 ;
        RECT 3.115 0.43 3.355 0.55 ;
        RECT 3.115 -0.18 3.235 0.55 ;
        RECT 2.275 -0.18 2.395 0.71 ;
        RECT 1.435 -0.18 1.555 0.71 ;
        RECT 0.535 -0.18 0.655 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 10.715 1.74 10.835 2.79 ;
        RECT 9.335 1.6 9.455 2.79 ;
        RECT 7.345 1.85 7.465 2.79 ;
        RECT 5.275 2.07 5.515 2.19 ;
        RECT 5.275 2.07 5.395 2.79 ;
        RECT 3.435 2.01 3.675 2.13 ;
        RECT 3.435 2.01 3.555 2.79 ;
        RECT 2.475 2.01 2.715 2.13 ;
        RECT 2.475 2.01 2.595 2.79 ;
        RECT 1.515 2.01 1.755 2.13 ;
        RECT 1.515 2.01 1.635 2.79 ;
        RECT 0.615 2.11 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.46 1.5 11.36 1.5 11.36 1.8 11.24 1.8 11.24 1.62 10.215 1.62 10.215 1.24 10.335 1.24 10.335 1.5 11.24 1.5 11.24 1.38 11.34 1.38 11.34 0.58 11.46 0.58 ;
      POLYGON 10.4 0.85 9.855 0.85 9.855 1.08 9.74 1.08 9.74 1.56 10.095 1.56 10.095 2.21 9.975 2.21 9.975 1.68 9.62 1.68 9.62 1.48 8.785 1.48 8.785 1.56 8.585 1.56 8.585 2.01 8.465 2.01 8.465 1.44 8.665 1.44 8.665 0.84 8.625 0.84 8.625 0.6 8.745 0.6 8.745 0.72 8.785 0.72 8.785 1.36 9.62 1.36 9.62 0.96 9.735 0.96 9.735 0.73 10.28 0.73 10.28 0.59 10.4 0.59 ;
      POLYGON 9.135 0.68 9.015 0.68 9.015 0.48 8.505 0.48 8.505 0.96 8.545 0.96 8.545 1.32 8.345 1.32 8.345 2.13 8.855 2.13 8.855 1.68 8.975 1.68 8.975 2.25 8.225 2.25 8.225 1.32 8.005 1.32 8.005 1.44 7.885 1.44 7.885 1.2 8.425 1.2 8.425 1.08 8.385 1.08 8.385 0.36 9.135 0.36 ;
      POLYGON 8.265 1.05 7.765 1.05 7.765 1.56 8.105 1.56 8.105 2.21 7.985 2.21 7.985 1.68 6.715 1.68 6.715 1.82 6.595 1.82 6.595 1.49 6.655 1.49 6.655 0.75 6.635 0.75 6.635 0.63 6.875 0.63 6.875 0.75 6.775 0.75 6.775 1.56 7.645 1.56 7.645 0.93 8.145 0.93 8.145 0.62 8.265 0.62 ;
      POLYGON 7.205 0.81 7.085 0.81 7.085 0.51 6.515 0.51 6.515 1.13 6.535 1.13 6.535 1.37 6.475 1.37 6.475 1.94 6.985 1.94 6.985 2.03 7.105 2.03 7.105 2.15 6.865 2.15 6.865 2.06 6.355 2.06 6.355 1.13 6.395 1.13 6.395 0.51 5.915 0.51 5.915 0.91 5.995 0.91 5.995 1.15 5.795 1.15 5.795 0.61 5.035 0.61 5.035 0.51 4.555 0.51 4.555 0.97 4.815 0.97 4.815 1.09 4.435 1.09 4.435 0.39 5.155 0.39 5.155 0.49 5.795 0.49 5.795 0.39 7.205 0.39 ;
      POLYGON 6.275 0.75 6.235 0.75 6.235 1.99 6.115 1.99 6.115 1.39 5.315 1.39 5.315 1.31 5.175 1.31 5.175 1.19 5.435 1.19 5.435 1.27 6.115 1.27 6.115 0.75 6.035 0.75 6.035 0.63 6.275 0.63 ;
      POLYGON 6.075 2.25 5.835 2.25 5.835 1.95 4.555 1.95 4.555 2.23 3.905 2.23 3.905 1.89 0.135 1.89 0.135 1.71 0.12 1.71 0.12 0.78 0.135 0.78 0.135 0.66 0.255 0.66 0.255 0.9 0.24 0.9 0.24 1.59 0.255 1.59 0.255 1.77 3.715 1.77 3.715 0.91 3.835 0.91 3.835 1.77 4.025 1.77 4.025 2.11 4.435 2.11 4.435 1.33 4.215 1.33 4.215 1.21 4.555 1.21 4.555 1.83 5.955 1.83 5.955 2.13 6.075 2.13 ;
      POLYGON 5.675 1.15 5.555 1.15 5.555 1.07 5.055 1.07 5.055 1.59 4.975 1.59 4.975 1.71 4.855 1.71 4.855 1.47 4.935 1.47 4.935 0.85 4.675 0.85 4.675 0.63 4.915 0.63 4.915 0.73 5.055 0.73 5.055 0.95 5.555 0.95 5.555 0.91 5.675 0.91 ;
      POLYGON 4.315 1.99 4.195 1.99 4.195 1.59 3.975 1.59 3.975 0.79 3.095 0.79 3.095 1.13 2.975 1.13 2.975 0.67 3.975 0.67 3.975 0.57 4.095 0.57 4.095 1.47 4.315 1.47 ;
      POLYGON 3.515 1.37 2.855 1.37 2.855 1.53 3.195 1.53 3.195 1.65 2.735 1.65 2.735 1.25 2.075 1.25 2.075 1.13 2.735 1.13 2.735 0.81 2.695 0.81 2.695 0.57 2.815 0.57 2.815 0.69 2.855 0.69 2.855 1.25 3.395 1.25 3.395 0.91 3.515 0.91 ;
  END
END SMDFFHQX4

MACRO BUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1 1.67 1.5 ;
        RECT 1.52 1 1.67 1.47 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.32 1.095 2.21 ;
        RECT 0.975 0.4 1.095 0.64 ;
        RECT 0.135 0.76 1.09 0.88 ;
        RECT 0.135 1.32 1.095 1.44 ;
        RECT 0.97 0.52 1.09 0.88 ;
        RECT 0.36 1.175 0.51 1.44 ;
        RECT 0.36 0.76 0.48 1.44 ;
        RECT 0.135 1.32 0.255 2.21 ;
        RECT 0.135 0.59 0.255 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.395 1.62 1.515 2.79 ;
        RECT 0.555 1.56 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 2.21 1.815 2.21 1.815 0.88 1.33 0.88 1.33 1.17 1.21 1.17 1.21 0.76 1.815 0.76 1.815 0.59 1.935 0.59 ;
  END
END BUFX3

MACRO AOI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.99 1.775 1.11 ;
        RECT 0.595 0.94 1.62 0.99 ;
        RECT 0.735 0.87 1.62 0.99 ;
        RECT 0.555 0.97 0.855 1.09 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 0.94 3.465 1.09 ;
        RECT 3.095 0.94 3.335 1.11 ;
        RECT 2.44 0.87 3.325 0.99 ;
        RECT 2.135 0.99 2.56 1.11 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.14 2.83 1.61 ;
        RECT 2.68 1.11 2.8 1.61 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.11 1.38 1.58 ;
        RECT 1.255 1.11 1.375 1.61 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 1.56 3.215 2.01 ;
        RECT 2.255 1.73 3.215 1.85 ;
        RECT 1.055 0.63 2.855 0.75 ;
        RECT 2.255 1.26 2.375 2.01 ;
        RECT 1.755 1.26 2.375 1.38 ;
        RECT 1.755 1.23 2.015 1.38 ;
        RECT 1.895 0.63 2.015 1.38 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.315 -0.18 3.435 0.64 ;
        RECT 1.835 0.39 2.075 0.51 ;
        RECT 1.835 -0.18 1.955 0.51 ;
        RECT 0.475 -0.18 0.595 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 1.415 1.97 1.535 2.79 ;
        RECT 0.575 1.97 0.695 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.635 2.25 1.835 2.25 1.835 1.85 1.115 1.85 1.115 2.21 0.995 2.21 0.995 1.85 0.275 1.85 0.275 2.21 0.155 2.21 0.155 1.56 0.275 1.56 0.275 1.73 0.995 1.73 0.995 1.7 1.115 1.7 1.115 1.73 1.835 1.73 1.835 1.56 1.955 1.56 1.955 2.13 2.675 2.13 2.675 1.97 2.795 1.97 2.795 2.13 3.515 2.13 3.515 1.56 3.635 1.56 ;
  END
END AOI22X2

MACRO MXI3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X4 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.255 1 0.375 1.24 ;
        RECT 0.07 1 0.375 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.285 1.41 2.565 1.53 ;
        RECT 2.285 1.09 2.405 1.53 ;
        RECT 1.725 1.09 2.405 1.21 ;
        RECT 1.805 0.885 1.96 1.21 ;
        RECT 1.725 1.09 1.845 1.34 ;
        RECT 1.245 1.18 1.925 1.3 ;
        RECT 1.125 1.3 1.365 1.42 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.685 1.2 4.805 1.44 ;
        RECT 4.42 1.2 4.805 1.435 ;
        RECT 4.42 1.175 4.57 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.965 1.23 6.365 1.48 ;
        RECT 6.105 1.21 6.365 1.48 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.345 0.97 6.525 1.09 ;
        RECT 5.725 0.94 6.075 1.09 ;
        RECT 5.725 0.93 5.845 1.17 ;
        RECT 5.165 1.38 5.465 1.5 ;
        RECT 5.345 0.97 5.465 1.5 ;
        RECT 5.165 1.38 5.285 1.62 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.445 0.69 4.645 0.81 ;
        RECT 4.185 1.555 4.305 2.21 ;
        RECT 4.18 0.69 4.3 1.675 ;
        RECT 3.525 1.32 4.3 1.44 ;
        RECT 3.55 1.175 3.7 1.44 ;
        RECT 3.345 1.46 3.645 1.58 ;
        RECT 3.525 1.32 3.645 1.58 ;
        RECT 3.345 1.46 3.465 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.285 -0.18 6.405 0.81 ;
        RECT 4.885 -0.18 5.125 0.33 ;
        RECT 3.925 -0.18 4.165 0.33 ;
        RECT 2.965 -0.18 3.085 0.68 ;
        RECT 1.465 -0.18 1.585 0.68 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 6.085 1.84 6.205 2.79 ;
        RECT 4.605 1.56 4.725 2.79 ;
        RECT 3.765 1.56 3.885 2.79 ;
        RECT 2.925 1.56 3.045 2.79 ;
        RECT 1.565 1.78 1.685 2.79 ;
        RECT 0.135 1.46 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.825 0.81 6.765 0.81 6.765 1.84 6.625 1.84 6.625 1.96 6.505 1.96 6.505 1.72 5.585 1.72 5.585 1.4 5.705 1.4 5.705 1.6 6.645 1.6 6.645 0.69 6.705 0.69 6.705 0.57 6.825 0.57 ;
      POLYGON 5.765 0.81 5.645 0.81 5.645 0.69 5.045 0.69 5.045 1.74 5.445 1.74 5.445 1.98 5.325 1.98 5.325 1.86 4.925 1.86 4.925 0.69 4.795 0.69 4.795 0.57 3.325 0.57 3.325 0.92 3.005 0.92 3.005 1.04 2.765 1.04 2.765 0.92 2.885 0.92 2.885 0.8 3.205 0.8 3.205 0.45 4.915 0.45 4.915 0.57 5.765 0.57 ;
      POLYGON 3.405 1.34 2.805 1.34 2.805 1.77 2.405 1.77 2.405 1.81 2.345 1.81 2.345 2.21 2.225 2.21 2.225 1.69 2.285 1.69 2.285 1.65 2.685 1.65 2.685 1.28 2.525 1.28 2.525 0.78 2.105 0.78 2.105 0.54 2.225 0.54 2.225 0.66 2.645 0.66 2.645 1.16 2.805 1.16 2.805 1.22 3.405 1.22 ;
      POLYGON 2.165 1.57 2.105 1.57 2.105 1.66 1.145 1.66 1.145 1.93 1.025 1.93 1.025 1.78 0.885 1.78 0.885 0.72 0.865 0.72 0.865 0.6 1.105 0.6 1.105 0.72 1.005 0.72 1.005 1.54 1.985 1.54 1.985 1.45 2.045 1.45 2.045 1.33 2.165 1.33 ;
      POLYGON 1.585 1.06 1.345 1.06 1.345 0.92 1.225 0.92 1.225 0.48 0.655 0.48 0.655 0.8 0.675 0.8 0.675 1.58 0.555 1.58 0.555 0.92 0.535 0.92 0.535 0.36 1.345 0.36 1.345 0.8 1.465 0.8 1.465 0.94 1.585 0.94 ;
  END
END MXI3X4

MACRO TLATNCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX2 0 0 ;
  SIZE 5.8 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 1.02 0.8 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
        RECT 0.445 1.02 0.565 1.26 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.655 1.23 4.915 1.45 ;
        RECT 4.655 1.18 4.775 1.57 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.095 1.145 1.215 1.58 ;
        RECT 0.94 0.885 1.185 1.145 ;
        RECT 1.065 0.68 1.185 1.265 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.8 0.18 ;
        RECT 4.735 0.46 4.975 0.58 ;
        RECT 4.735 -0.18 4.855 0.58 ;
        RECT 3.055 -0.18 3.175 0.38 ;
        RECT 1.485 -0.18 1.605 0.73 ;
        RECT 0.645 -0.18 0.765 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.8 2.79 ;
        RECT 4.735 1.69 4.855 2.79 ;
        RECT 3.255 2.11 3.375 2.79 ;
        RECT 2.295 2.12 2.415 2.79 ;
        RECT 1.515 2.12 1.755 2.24 ;
        RECT 1.515 2.12 1.635 2.79 ;
        RECT 0.615 1.94 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.395 1.75 5.095 1.75 5.095 1.63 5.275 1.63 5.275 0.82 4.495 0.82 4.495 0.52 3.335 0.52 3.335 0.4 4.615 0.4 4.615 0.7 5.275 0.7 5.275 0.66 5.395 0.66 ;
      POLYGON 5.155 1.24 5.035 1.24 5.035 1.06 4.535 1.06 4.535 1.71 4.275 1.71 4.275 1.75 4.035 1.75 4.035 1.63 4.155 1.63 4.155 1.59 4.415 1.59 4.415 1.06 3.895 1.06 3.895 0.66 4.015 0.66 4.015 0.94 5.155 0.94 ;
      POLYGON 4.295 1.47 4.175 1.47 4.175 1.35 2.165 1.35 2.165 1.52 1.925 1.52 1.925 1.4 1.965 1.4 1.965 0.68 2.085 0.68 2.085 1.23 3.635 1.23 3.635 1 3.755 1 3.755 1.23 4.295 1.23 ;
      POLYGON 3.935 2.25 3.815 2.25 3.815 1.99 2.875 1.99 2.875 2 1.04 2 1.04 1.82 0.135 1.82 0.135 1.46 0.165 1.46 0.165 0.68 0.285 0.68 0.285 1.58 0.255 1.58 0.255 1.7 1.16 1.7 1.16 1.88 2.755 1.88 2.755 1.87 3.935 1.87 ;
      POLYGON 2.955 1.75 2.57 1.75 2.57 1.76 1.685 1.76 1.685 1.2 1.335 1.2 1.335 1.08 1.685 1.08 1.685 0.85 1.725 0.85 1.725 0.44 2.475 0.44 2.475 0.9 2.355 0.9 2.355 0.56 1.845 0.56 1.845 0.97 1.805 0.97 1.805 1.64 2.45 1.64 2.45 1.63 2.955 1.63 ;
  END
END TLATNCAX2

MACRO OAI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X2 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.175 2.83 1.435 ;
        RECT 2.515 1.175 2.83 1.295 ;
        RECT 2.515 1.055 2.635 1.295 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1 2.155 1.15 ;
        RECT 1.755 0.94 2.015 1.12 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 1.04 1.635 1.16 ;
        RECT 0.65 1.04 0.8 1.435 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.555 1.515 2.21 ;
        RECT 0.07 1.555 1.515 1.675 ;
        RECT 0.195 0.8 1.095 0.92 ;
        RECT 0.975 0.63 1.095 0.92 ;
        RECT 0.555 1.555 0.675 2.21 ;
        RECT 0.195 0.8 0.315 1.675 ;
        RECT 0.07 1.465 0.22 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.615 -0.18 1.735 0.68 ;
        RECT 0.335 -0.18 0.455 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.645 2.2 2.765 2.79 ;
        RECT 1.875 2.2 1.995 2.79 ;
        RECT 0.975 1.795 1.095 2.79 ;
        RECT 0.135 1.845 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.635 0.81 2.395 0.81 2.395 1.52 2.355 1.52 2.355 1.8 2.235 1.8 2.235 1.4 1.075 1.4 1.075 1.28 2.275 1.28 2.275 0.69 2.635 0.69 ;
  END
END OAI2BB1X2

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 1.26 1.4 1.38 ;
        RECT 0.885 1.23 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.52 0.85 1.64 1.725 ;
        RECT 1.5 1.5 1.62 2.21 ;
        RECT 0.66 0.85 1.64 0.97 ;
        RECT 1.5 0.68 1.62 0.97 ;
        RECT 0.66 1.5 1.67 1.62 ;
        RECT 0.66 1.5 0.78 2.21 ;
        RECT 0.66 0.68 0.78 0.97 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.92 -0.18 2.04 0.73 ;
        RECT 1.08 -0.18 1.2 0.73 ;
        RECT 0.24 -0.18 0.36 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.92 1.56 2.04 2.79 ;
        RECT 1.08 1.74 1.2 2.79 ;
        RECT 0.24 1.56 0.36 2.79 ;
    END
  END VDD
END INVX4

MACRO FILL64
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL64 0 0 ;
  SIZE 18.56 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 18.56 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 18.56 0.18 ;
    END
  END VSS
END FILL64

MACRO TLATNCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX20 0 0 ;
  SIZE 15.37 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.06 0.51 1.525 ;
        RECT 0.38 1.03 0.5 1.525 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.135 0.84 1.525 ;
        RECT 0.72 1.12 0.84 1.525 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6387 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.09 1.205 15.21 2.205 ;
        RECT 15.01 0.405 15.13 1.03 ;
        RECT 8.19 1.205 15.21 1.325 ;
        RECT 14.83 0.91 15.13 1.03 ;
        RECT 14.17 1.03 14.95 1.325 ;
        RECT 14.25 1.03 14.37 2.21 ;
        RECT 14.17 0.405 14.29 1.325 ;
        RECT 13.41 1.205 13.53 2.21 ;
        RECT 13.15 0.79 13.45 0.91 ;
        RECT 13.33 0.405 13.45 0.91 ;
        RECT 12.49 1.03 13.27 1.325 ;
        RECT 13.15 0.79 13.27 1.325 ;
        RECT 12.57 1.03 12.69 2.21 ;
        RECT 12.49 0.405 12.61 1.325 ;
        RECT 11.73 1.205 11.85 2.21 ;
        RECT 11.47 0.79 11.77 0.91 ;
        RECT 11.65 0.405 11.77 0.91 ;
        RECT 10.81 1.03 11.59 1.325 ;
        RECT 11.47 0.79 11.59 1.325 ;
        RECT 10.89 1.03 11.01 2.21 ;
        RECT 10.81 0.405 10.93 1.325 ;
        RECT 10.05 1.205 10.17 2.21 ;
        RECT 9.79 0.79 10.09 0.91 ;
        RECT 9.97 0.405 10.09 0.91 ;
        RECT 9.07 1.03 9.91 1.325 ;
        RECT 9.79 0.79 9.91 1.325 ;
        RECT 9.21 1.03 9.33 2.21 ;
        RECT 9.07 0.4 9.19 1.325 ;
        RECT 8.37 1.205 8.49 2.21 ;
        RECT 8.23 1.205 8.49 1.445 ;
        RECT 8.19 1.175 8.35 1.435 ;
        RECT 8.23 0.4 8.35 1.445 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 15.37 0.18 ;
        RECT 14.59 -0.18 14.71 0.91 ;
        RECT 13.75 -0.18 13.87 0.91 ;
        RECT 12.91 -0.18 13.03 0.91 ;
        RECT 12.07 -0.18 12.19 0.91 ;
        RECT 11.23 -0.18 11.35 0.91 ;
        RECT 10.39 -0.18 10.51 0.91 ;
        RECT 9.55 -0.18 9.67 0.91 ;
        RECT 8.65 -0.18 8.77 0.91 ;
        RECT 7.81 -0.18 7.93 0.87 ;
        RECT 6.21 0.46 6.45 0.58 ;
        RECT 6.21 -0.18 6.33 0.58 ;
        RECT 4.73 0.46 4.97 0.58 ;
        RECT 4.73 -0.18 4.85 0.58 ;
        RECT 2.975 -0.18 3.215 0.32 ;
        RECT 2.015 -0.18 2.255 0.32 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 15.37 2.79 ;
        RECT 14.67 1.445 14.79 2.79 ;
        RECT 13.83 1.445 13.95 2.79 ;
        RECT 12.99 1.445 13.11 2.79 ;
        RECT 12.15 1.445 12.27 2.79 ;
        RECT 11.31 1.445 11.43 2.79 ;
        RECT 10.47 1.445 10.59 2.79 ;
        RECT 9.63 1.445 9.75 2.79 ;
        RECT 8.79 1.445 8.91 2.79 ;
        RECT 7.95 1.71 8.07 2.79 ;
        RECT 7.11 1.71 7.23 2.79 ;
        RECT 6.27 1.71 6.39 2.79 ;
        RECT 5.43 1.71 5.55 2.79 ;
        RECT 4.59 1.71 4.71 2.79 ;
        RECT 3.75 1.91 3.87 2.79 ;
        RECT 2.9 2.15 3.14 2.27 ;
        RECT 2.9 2.15 3.02 2.79 ;
        RECT 1.94 1.97 2.18 2.09 ;
        RECT 1.94 1.97 2.06 2.79 ;
        RECT 0.66 1.645 0.78 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.07 1.23 8.01 1.23 8.01 1.59 7.65 1.59 7.65 2.21 7.53 2.21 7.53 1.59 6.81 1.59 6.81 2.21 6.69 2.21 6.69 1.59 5.97 1.59 5.97 2.21 5.85 2.21 5.85 1.59 5.13 1.59 5.13 2.21 5.01 2.21 5.01 1.59 4.29 1.59 4.29 2.21 4.17 2.21 4.17 1.47 7.89 1.47 7.89 1.11 7.15 1.11 7.15 0.83 7.11 0.83 7.11 0.82 4.21 0.82 4.21 0.77 4.09 0.77 4.09 0.65 4.33 0.65 4.33 0.7 5.37 0.7 5.37 0.65 5.61 0.65 5.61 0.7 7.11 0.7 7.11 0.59 7.23 0.59 7.23 0.71 7.27 0.71 7.27 0.99 8.07 0.99 ;
      POLYGON 7.77 1.35 4.05 1.35 4.05 1.79 3.01 1.79 3.01 1.61 2.48 1.61 2.48 1.37 2.595 1.37 2.595 0.95 1.795 0.95 1.795 0.83 2.495 0.83 2.495 0.68 2.735 0.68 2.735 0.8 2.715 0.8 2.715 1.49 3.13 1.49 3.13 1.67 3.93 1.67 3.93 1.23 7.77 1.23 ;
      POLYGON 7.03 1.11 3.635 1.11 3.635 1.55 3.38 1.55 3.38 1.43 3.515 1.43 3.515 0.56 1.655 0.56 1.655 1.01 1.535 1.01 1.535 0.44 3.635 0.44 3.635 0.99 7.03 0.99 ;
      POLYGON 3.46 2.03 2.645 2.03 2.645 1.85 1.705 1.85 1.705 2.005 1.58 2.005 1.58 2.225 1.46 2.225 1.46 2.005 1.055 2.005 1.055 0.91 0.24 0.91 0.24 1.645 0.36 1.645 0.36 1.885 0.24 1.885 0.24 1.765 0.12 1.765 0.12 0.67 0.135 0.67 0.135 0.43 0.255 0.43 0.255 0.79 1.055 0.79 1.055 0.75 1.175 0.75 1.175 1.885 1.585 1.885 1.585 1.73 2.765 1.73 2.765 1.91 3.46 1.91 ;
      POLYGON 2.475 1.25 1.42 1.25 1.42 1.765 1.3 1.765 1.3 1.37 1.295 1.37 1.295 0.43 1.415 0.43 1.415 1.13 2.235 1.13 2.235 1.09 2.475 1.09 ;
  END
END TLATNCAX20

MACRO INVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX20 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.16 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.165 6.365 1.285 ;
        RECT 0.885 1.165 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.285 1.45 7.405 2.21 ;
        RECT 0.555 0.925 7.405 1.045 ;
        RECT 7.285 0.4 7.405 1.045 ;
        RECT 0.565 1.5 7.405 1.62 ;
        RECT 6.74 1.175 6.89 1.62 ;
        RECT 6.485 1.315 6.89 1.62 ;
        RECT 6.485 0.925 6.605 1.62 ;
        RECT 6.445 1.445 6.565 2.21 ;
        RECT 6.445 0.4 6.565 1.045 ;
        RECT 5.605 1.445 5.725 2.21 ;
        RECT 5.605 0.4 5.725 1.045 ;
        RECT 4.765 1.445 4.885 2.21 ;
        RECT 4.765 0.4 4.885 1.045 ;
        RECT 3.925 1.445 4.045 2.21 ;
        RECT 3.925 0.4 4.045 1.045 ;
        RECT 3.085 1.445 3.205 2.21 ;
        RECT 3.085 0.4 3.205 1.045 ;
        RECT 2.245 1.445 2.365 2.21 ;
        RECT 2.245 0.4 2.365 1.045 ;
        RECT 1.405 1.445 1.525 2.21 ;
        RECT 1.395 0.4 1.515 1.045 ;
        RECT 0.565 1.445 0.685 2.21 ;
        RECT 0.555 0.4 0.675 1.045 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.865 -0.18 6.985 0.805 ;
        RECT 6.025 -0.18 6.145 0.805 ;
        RECT 5.185 -0.18 5.305 0.805 ;
        RECT 4.345 -0.18 4.465 0.805 ;
        RECT 3.505 -0.18 3.625 0.805 ;
        RECT 2.665 -0.18 2.785 0.805 ;
        RECT 1.825 -0.18 1.945 0.805 ;
        RECT 0.975 -0.18 1.095 0.805 ;
        RECT 0.135 -0.18 0.255 0.91 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.865 1.74 6.985 2.79 ;
        RECT 6.025 1.74 6.145 2.79 ;
        RECT 5.185 1.74 5.305 2.79 ;
        RECT 4.345 1.74 4.465 2.79 ;
        RECT 3.505 1.74 3.625 2.79 ;
        RECT 2.665 1.74 2.785 2.79 ;
        RECT 1.825 1.74 1.945 2.79 ;
        RECT 0.985 1.74 1.105 2.79 ;
        RECT 0.145 1.445 0.265 2.79 ;
    END
  END VDD
END INVX20

MACRO AOI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.525 0.99 8.525 1.11 ;
        RECT 5.525 0.94 5.785 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.925 0.99 5.165 1.11 ;
        RECT 5 0.885 5.15 1.145 ;
        RECT 5 0.75 5.12 1.145 ;
        RECT 0.745 0.75 5.12 0.87 ;
        RECT 2.905 0.75 3.145 1.09 ;
        RECT 0.745 0.75 0.865 1.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 1 4.805 1.12 ;
        RECT 2.665 1.21 3.58 1.33 ;
        RECT 3.46 1 3.58 1.33 ;
        RECT 2.665 1.06 2.785 1.33 ;
        RECT 2.135 1.06 2.785 1.18 ;
        RECT 1.025 0.99 2.255 1.11 ;
        RECT 1.23 0.99 1.38 1.435 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.185 1.26 7.785 1.38 ;
        RECT 6.395 1.23 6.655 1.38 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.425 1.45 3.925 1.57 ;
        RECT 3.805 1.24 3.925 1.57 ;
        RECT 2.425 1.3 2.545 1.57 ;
        RECT 1.785 1.3 2.545 1.42 ;
        RECT 1.755 1.23 2.015 1.38 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.285 1.5 8.405 2.01 ;
        RECT 5.765 1.5 8.405 1.62 ;
        RECT 1.705 0.51 7.665 0.63 ;
        RECT 7.445 1.5 7.565 2.01 ;
        RECT 6.605 1.5 6.725 2.01 ;
        RECT 5.765 1.32 5.885 2.01 ;
        RECT 5.285 1.23 5.785 1.44 ;
        RECT 5.285 0.51 5.405 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.125 -0.18 8.245 0.64 ;
        RECT 6.725 -0.18 6.965 0.39 ;
        RECT 5.245 -0.18 5.485 0.39 ;
        RECT 2.725 -0.18 2.965 0.39 ;
        RECT 0.545 0.46 0.785 0.58 ;
        RECT 0.545 -0.18 0.665 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 4.925 1.93 5.045 2.79 ;
        RECT 4.085 1.93 4.205 2.79 ;
        RECT 3.245 1.93 3.365 2.79 ;
        RECT 2.405 1.93 2.525 2.79 ;
        RECT 1.565 1.93 1.685 2.79 ;
        RECT 0.725 1.93 0.845 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.825 2.25 5.345 2.25 5.345 1.81 4.625 1.81 4.625 2.21 4.505 2.21 4.505 1.81 3.785 1.81 3.785 2.21 3.665 2.21 3.665 1.81 2.945 1.81 2.945 2.21 2.825 2.21 2.825 1.81 2.105 1.81 2.105 2.21 1.985 2.21 1.985 1.81 1.265 1.81 1.265 2.21 1.145 2.21 1.145 1.81 0.425 1.81 0.425 2.21 0.305 2.21 0.305 1.56 0.425 1.56 0.425 1.69 1.145 1.69 1.145 1.56 1.265 1.56 1.265 1.69 1.985 1.69 1.985 1.56 2.105 1.56 2.105 1.69 4.505 1.69 4.505 1.56 4.625 1.56 4.625 1.69 5.345 1.69 5.345 1.56 5.465 1.56 5.465 2.13 6.185 2.13 6.185 1.74 6.305 1.74 6.305 2.13 7.025 2.13 7.025 1.74 7.145 1.74 7.145 2.13 7.865 2.13 7.865 1.74 7.985 1.74 7.985 2.13 8.705 2.13 8.705 1.56 8.825 1.56 ;
  END
END AOI32X4

MACRO SDFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX1 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.22 0.895 1.46 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.34 0.8 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.605 1.21 5.725 1.45 ;
        RECT 5.235 1.23 5.725 1.38 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.685 1.21 7.045 1.41 ;
        RECT 6.685 1.21 6.945 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.205 0.89 7.345 1.01 ;
        RECT 6.975 0.89 7.235 1.09 ;
        RECT 6.505 0.77 6.625 1.01 ;
        RECT 6.205 0.89 6.325 1.43 ;
        RECT 6.085 1.31 6.205 1.55 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 2.21 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.005 1.97 7.125 2.79 ;
        RECT 5.725 1.97 5.845 2.79 ;
        RECT 3.675 2.2 3.795 2.79 ;
        RECT 2.015 2.14 2.255 2.26 ;
        RECT 2.015 2.14 2.135 2.79 ;
        RECT 0.555 1.845 0.675 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.005 -0.18 7.125 0.65 ;
        RECT 5.725 -0.18 5.845 0.65 ;
        RECT 3.615 -0.18 3.855 0.34 ;
        RECT 1.875 -0.18 2.115 0.32 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.585 1.795 7.545 1.795 7.545 2.09 7.425 2.09 7.425 1.675 6.445 1.675 6.445 1.13 6.565 1.13 6.565 1.555 7.465 1.555 7.465 0.77 7.425 0.77 7.425 0.41 7.545 0.41 7.545 0.65 7.585 0.65 ;
      POLYGON 6.485 0.65 6.085 0.65 6.085 1.19 5.965 1.19 5.965 1.67 6.325 1.67 6.325 1.795 6.485 1.795 6.485 2.09 6.365 2.09 6.365 1.915 6.205 1.915 6.205 1.79 4.855 1.79 4.855 1.67 4.915 1.67 4.915 0.68 5.035 0.68 5.035 1.67 5.845 1.67 5.845 1.07 5.965 1.07 5.965 0.53 6.365 0.53 6.365 0.41 6.485 0.41 ;
      POLYGON 5.485 2.03 4.615 2.03 4.615 1.28 4.675 1.28 4.675 0.56 4.175 0.56 4.175 0.58 3.115 0.58 3.115 1.24 2.995 1.24 2.995 0.46 4.055 0.46 4.055 0.44 4.155 0.44 4.155 0.4 4.395 0.4 4.395 0.44 5.305 0.44 5.305 0.41 5.425 0.41 5.425 0.65 5.305 0.65 5.305 0.56 4.795 0.56 4.795 1.52 4.735 1.52 4.735 1.91 5.485 1.91 ;
      POLYGON 4.555 0.86 4.495 0.86 4.495 1.84 4.375 1.84 4.375 1.44 3.495 1.44 3.495 1.32 4.375 1.32 4.375 0.86 4.315 0.86 4.315 0.74 4.555 0.74 ;
      POLYGON 4.415 2.22 3.985 2.22 3.985 2.08 3.165 2.08 3.165 2.22 2.925 2.22 2.925 2.08 2.395 2.08 2.395 2.02 1.035 2.02 1.035 0.68 1.155 0.68 1.155 1.9 2.395 1.9 2.395 1.06 2.635 1.06 2.635 1.18 2.515 1.18 2.515 1.96 4.105 1.96 4.105 2.1 4.415 2.1 ;
      POLYGON 4.075 1.2 3.355 1.2 3.355 1.72 3.315 1.72 3.315 1.84 3.195 1.84 3.195 1.6 3.235 1.6 3.235 0.74 3.475 0.74 3.475 0.86 3.355 0.86 3.355 1.08 4.075 1.08 ;
      POLYGON 2.895 1.84 2.775 1.84 2.775 1.48 2.755 1.48 2.755 0.92 2.715 0.92 2.715 0.68 1.665 0.68 1.665 0.56 1.515 0.56 1.515 0.4 1.755 0.4 1.755 0.44 1.785 0.44 1.785 0.56 2.835 0.56 2.835 0.8 2.875 0.8 2.875 1.36 2.895 1.36 ;
      POLYGON 2.275 1.26 1.655 1.26 1.655 1.66 1.775 1.66 1.775 1.78 1.535 1.78 1.535 0.92 1.425 0.92 1.425 0.8 1.275 0.8 1.275 0.56 0.915 0.56 0.915 1.1 0.535 1.1 0.535 1.24 0.415 1.24 0.415 0.98 0.795 0.98 0.795 0.44 1.395 0.44 1.395 0.68 1.545 0.68 1.545 0.8 1.655 0.8 1.655 1.14 2.275 1.14 ;
  END
END SDFFQX1

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.935 1.36 ;
        RECT 0.815 1.12 0.935 1.36 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.615 1.26 2.855 1.38 ;
        RECT 1.955 1.28 2.735 1.4 ;
        RECT 2.045 1.23 2.305 1.4 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.885 0.455 1.025 ;
        RECT 0.335 0.68 0.455 1.025 ;
        RECT 0.135 0.885 0.255 2.19 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.455 0.68 2.695 0.8 ;
        RECT 2.535 -0.18 2.655 0.8 ;
        RECT 0.755 -0.18 0.875 0.86 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.395 2.24 2.635 2.79 ;
        RECT 0.615 2.18 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.095 1.66 3.055 1.66 3.055 1.9 1.995 1.9 1.995 2.2 1.175 2.2 1.175 2.08 1.875 2.08 1.875 1.78 2.935 1.78 2.935 1.54 2.975 1.54 2.975 1.11 1.795 1.11 1.795 1.22 1.675 1.22 1.675 0.98 1.795 0.98 1.795 0.99 2.935 0.99 2.935 0.62 3.055 0.62 3.055 0.87 3.095 0.87 ;
      POLYGON 2.415 0.48 1.295 0.48 1.295 1.72 0.915 1.72 0.915 1.6 1.175 1.6 1.175 0.36 2.415 0.36 ;
      POLYGON 1.715 0.86 1.535 0.86 1.535 1.96 0.675 1.96 0.675 1.675 0.41 1.675 0.41 1.22 0.53 1.22 0.53 1.555 0.795 1.555 0.795 1.84 1.415 1.84 1.415 0.74 1.595 0.74 1.595 0.62 1.715 0.62 ;
  END
END XNOR2X1

MACRO CLKMX2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X12 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.194 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 1.415 1.27 1.535 ;
        RECT 0.39 1.555 1.11 1.675 ;
        RECT 0.99 1.415 1.11 1.675 ;
        RECT 0.39 1.175 0.51 1.675 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.095 0.87 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.93 1.215 2.25 1.435 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.93 1.215 2.05 1.455 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 1.31 6.07 2.21 ;
        RECT 5.77 1.31 6.07 1.43 ;
        RECT 5.79 0.405 5.91 1.16 ;
        RECT 2.61 1.19 5.89 1.31 ;
        RECT 4.95 1.04 5.89 1.31 ;
        RECT 5.11 1.04 5.23 2.21 ;
        RECT 4.95 0.405 5.07 1.31 ;
        RECT 4.27 1.19 4.39 2.21 ;
        RECT 3.27 1.04 4.23 1.31 ;
        RECT 4.11 0.405 4.23 1.31 ;
        RECT 3.43 1.04 3.55 2.21 ;
        RECT 3.27 0.405 3.39 1.31 ;
        RECT 2.61 1.175 2.83 1.435 ;
        RECT 2.61 0.695 2.73 1.48 ;
        RECT 2.59 1.36 2.71 2.21 ;
        RECT 2.37 0.46 2.61 0.815 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 6.21 -0.18 6.33 0.92 ;
        RECT 5.37 -0.18 5.49 0.92 ;
        RECT 4.53 -0.18 4.65 0.92 ;
        RECT 3.69 -0.18 3.81 0.92 ;
        RECT 2.85 -0.18 2.97 0.92 ;
        RECT 1.95 0.46 2.19 0.815 ;
        RECT 1.95 -0.18 2.07 0.815 ;
        RECT 0.61 -0.18 0.73 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 6.37 1.43 6.49 2.79 ;
        RECT 5.53 1.43 5.65 2.79 ;
        RECT 4.69 1.43 4.81 2.79 ;
        RECT 3.85 1.43 3.97 2.79 ;
        RECT 3.01 1.43 3.13 2.79 ;
        RECT 2.17 1.555 2.29 2.79 ;
        RECT 0.59 1.795 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.49 1.24 2.37 1.24 2.37 1.055 1.81 1.055 1.81 1.84 1.43 1.84 1.43 2.21 1.31 2.21 1.31 1.72 1.69 1.72 1.69 1.055 1.41 1.055 1.41 0.735 1.25 0.735 1.25 0.495 1.37 0.495 1.37 0.615 1.53 0.615 1.53 0.935 2.49 0.935 ;
      POLYGON 1.57 1.6 1.45 1.6 1.45 1.295 1.17 1.295 1.17 1 1.05 1 1.05 0.975 0.24 0.975 0.24 1.795 0.29 1.795 0.29 2.21 0.17 2.21 0.17 1.915 0.12 1.915 0.12 0.735 0.19 0.735 0.19 0.59 0.31 0.59 0.31 0.855 1.29 0.855 1.29 1.175 1.57 1.175 ;
  END
END CLKMX2X12

MACRO DFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRXL 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.875 1.48 2.115 1.64 ;
        RECT 1.755 1.52 2.015 1.715 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.59 1.23 7.65 1.35 ;
        RECT 6.05 1.12 6.71 1.24 ;
        RECT 6.05 0.4 6.17 1.24 ;
        RECT 5.085 0.4 6.17 0.52 ;
        RECT 3.28 1.16 5.205 1.28 ;
        RECT 5.085 0.4 5.205 1.28 ;
        RECT 4.945 0.94 5.205 1.28 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.35 1.12 9.555 1.435 ;
        RECT 9.35 1.07 9.525 1.435 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 1.04 10.66 1.45 ;
        RECT 10.525 1.04 10.645 1.525 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 0.92 ;
        RECT 1.355 1.32 1.475 2.09 ;
        RECT 1.335 0.8 1.455 1.44 ;
        RECT 1.23 0.885 1.455 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.705 -0.18 10.825 0.92 ;
        RECT 9.45 -0.18 9.57 0.89 ;
        RECT 7.75 -0.18 7.99 0.32 ;
        RECT 3.075 -0.18 3.195 0.78 ;
        RECT 1.785 -0.18 1.905 0.92 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.765 1.57 10.885 2.79 ;
        RECT 9.59 2.17 9.71 2.79 ;
        RECT 8.05 2.29 8.29 2.79 ;
        RECT 6.57 2.29 6.81 2.79 ;
        RECT 4.26 1.88 4.38 2.79 ;
        RECT 2.88 2.28 3.12 2.79 ;
        RECT 1.775 1.97 1.895 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.405 0.92 10.39 0.92 10.39 1.57 10.405 1.57 10.405 2.035 10.11 2.035 10.11 2.13 9.87 2.13 9.87 2.05 9.47 2.05 9.47 2.17 6.465 2.17 6.465 2.12 5.55 2.12 5.55 2 6.585 2 6.585 2.05 9.35 2.05 9.35 1.93 9.87 1.93 9.87 1.915 10.285 1.915 10.285 1.69 10.27 1.69 10.27 0.8 10.285 0.8 10.285 0.68 10.405 0.68 ;
      POLYGON 10.015 1.795 9.895 1.795 9.895 1.675 9.23 1.675 9.23 1.93 6.78 1.93 6.78 1.88 5.43 1.88 5.43 2.08 4.87 2.08 4.87 1.96 5.31 1.96 5.31 1.76 5.565 1.76 5.565 1.08 5.57 1.08 5.57 0.96 5.69 0.96 5.69 1.2 5.685 1.2 5.685 1.76 6.9 1.76 6.9 1.81 8.37 1.81 8.37 0.97 8.49 0.97 8.49 1.81 9.11 1.81 9.11 1.45 8.95 1.45 8.95 1.19 9.07 1.19 9.07 1.33 9.23 1.33 9.23 1.555 9.87 1.555 9.87 0.65 9.99 0.65 9.99 1.555 10.015 1.555 ;
      POLYGON 8.99 1.69 8.61 1.69 8.61 0.65 7.63 0.65 7.63 0.6 7.31 0.6 7.31 0.52 7.19 0.52 7.19 0.4 7.43 0.4 7.43 0.48 7.75 0.48 7.75 0.53 8.73 0.53 8.73 1.57 8.99 1.57 ;
      POLYGON 8.15 1.23 8.03 1.23 8.03 1.11 7.89 1.11 7.89 1.59 7.51 1.59 7.51 1.69 7.27 1.69 7.27 1.59 6.045 1.59 6.045 1.64 5.805 1.64 5.805 1.52 5.81 1.52 5.81 0.64 5.93 0.64 5.93 1.47 7.77 1.47 7.77 1.11 6.83 1.11 6.83 1 6.71 1 6.71 0.66 6.83 0.66 6.83 0.88 6.95 0.88 6.95 0.99 8.15 0.99 ;
      POLYGON 7.51 0.84 7.07 0.84 7.07 0.76 6.95 0.76 6.95 0.54 6.41 0.54 6.41 0.9 6.29 0.9 6.29 0.42 7.07 0.42 7.07 0.64 7.19 0.64 7.19 0.72 7.51 0.72 ;
      POLYGON 5.45 0.88 5.445 0.88 5.445 1.58 5.19 1.58 5.19 1.7 5.07 1.7 5.07 1.52 2.92 1.52 2.92 1.26 3.04 1.26 3.04 1.4 5.325 1.4 5.325 0.76 5.33 0.76 5.33 0.64 5.45 0.64 ;
      POLYGON 4.965 0.82 4.755 0.82 4.755 0.96 4.035 0.96 4.035 0.72 3.855 0.72 3.855 0.6 4.155 0.6 4.155 0.84 4.635 0.84 4.635 0.7 4.965 0.7 ;
      POLYGON 4.83 1.76 4.13 1.76 4.13 1.81 3.36 1.81 3.36 1.69 4.01 1.69 4.01 1.64 4.83 1.64 ;
      POLYGON 4.515 0.72 4.275 0.72 4.275 0.48 3.735 0.48 3.735 0.54 3.615 0.54 3.615 0.78 3.495 0.78 3.495 0.42 3.615 0.42 3.615 0.36 4.395 0.36 4.395 0.6 4.515 0.6 ;
      POLYGON 4.1 2.25 3.33 2.25 3.33 2.16 2.315 2.16 2.315 2.21 2.195 2.21 2.195 1.97 2.265 1.97 2.265 0.68 2.385 0.68 2.385 2.04 3.45 2.04 3.45 2.13 4.1 2.13 ;
      POLYGON 3.88 1.04 2.775 1.04 2.775 1.7 2.625 1.7 2.625 1.82 2.505 1.82 2.505 1.58 2.655 1.58 2.655 0.56 2.145 0.56 2.145 1.2 1.575 1.2 1.575 1.08 2.025 1.08 2.025 0.44 2.775 0.44 2.775 0.92 3.88 0.92 ;
      POLYGON 1.215 1.58 1.095 1.58 1.095 1.46 0.975 1.46 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 1.095 1.34 1.215 1.34 ;
  END
END DFFSRXL

MACRO DLY1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X4 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.15 0.565 1.38 ;
        RECT 0.305 1.15 0.425 1.56 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.385 1.36 3.505 2.13 ;
        RECT 2.68 0.76 3.505 0.88 ;
        RECT 3.385 0.59 3.505 0.88 ;
        RECT 3.205 1.36 3.505 1.48 ;
        RECT 2.68 1.24 3.325 1.36 ;
        RECT 2.68 1.175 2.83 1.435 ;
        RECT 2.545 1.36 2.8 1.48 ;
        RECT 2.68 0.71 2.8 1.48 ;
        RECT 2.545 0.71 2.8 0.83 ;
        RECT 2.545 1.36 2.665 2.13 ;
        RECT 2.545 0.59 2.665 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.805 -0.18 3.925 0.64 ;
        RECT 2.965 -0.18 3.085 0.64 ;
        RECT 2.125 -0.18 2.245 0.64 ;
        RECT 1.185 1.36 1.345 1.6 ;
        RECT 1.225 0.76 1.345 1.6 ;
        RECT 0.955 0.76 1.345 0.88 ;
        RECT 0.955 -0.18 1.075 0.88 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 3.805 1.48 3.925 2.79 ;
        RECT 2.965 1.48 3.085 2.79 ;
        RECT 2.125 1.48 2.245 2.79 ;
        RECT 0.985 1 1.105 1.24 ;
        RECT 0.945 1.12 1.065 2.79 ;
        RECT 0.555 1.82 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.385 1.15 2.285 1.15 2.285 1.36 1.825 1.36 1.825 2.13 1.705 2.13 1.705 1.24 2.165 1.24 2.165 0.88 1.705 0.88 1.705 0.59 1.825 0.59 1.825 0.76 2.385 0.76 ;
      POLYGON 2.045 1.12 1.585 1.12 1.585 1.84 1.315 1.84 1.315 1.96 1.195 1.96 1.195 1.72 1.465 1.72 1.465 0.64 1.195 0.64 1.195 0.4 1.315 0.4 1.315 0.52 1.585 0.52 1.585 1 2.045 1 ;
      POLYGON 0.825 1.03 0.185 1.03 0.185 1.68 0.255 1.68 0.255 1.94 0.135 1.94 0.135 1.8 0.065 1.8 0.065 0.52 0.135 0.52 0.135 0.4 0.255 0.4 0.255 0.64 0.185 0.64 0.185 0.91 0.825 0.91 ;
  END
END DLY1X4

MACRO MXI3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X2 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.395 1.295 ;
        RECT 0.275 1.055 0.395 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.52 2.95 1.64 ;
        RECT 2.83 1.24 2.95 1.64 ;
        RECT 2.29 1.02 2.41 1.64 ;
        RECT 2.045 1.52 2.305 1.67 ;
        RECT 1.23 1.26 1.35 1.64 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.13 1.175 4.53 1.295 ;
        RECT 4.41 1.055 4.53 1.295 ;
        RECT 4.13 1.175 4.28 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.87 1.11 6.05 1.5 ;
        RECT 5.93 1.1 6.05 1.5 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.395 0.94 6.655 1.09 ;
        RECT 5.11 0.86 6.515 0.98 ;
        RECT 6.29 0.94 6.655 1.06 ;
        RECT 5.61 0.84 5.73 1.08 ;
        RECT 4.89 1.4 5.23 1.52 ;
        RECT 5.11 0.86 5.23 1.52 ;
        RECT 4.89 1.4 5.01 1.64 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.81 0.74 4.05 0.86 ;
        RECT 3.87 0.74 3.99 2.21 ;
        RECT 3.84 1.175 3.99 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.09 -0.18 6.21 0.74 ;
        RECT 4.29 -0.18 4.53 0.38 ;
        RECT 3.33 -0.18 3.57 0.38 ;
        RECT 1.43 -0.18 1.55 0.38 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 5.99 1.86 6.11 2.79 ;
        RECT 4.29 1.56 4.41 2.79 ;
        RECT 3.45 1.58 3.57 2.79 ;
        RECT 1.43 2.22 1.55 2.79 ;
        RECT 0.135 1.555 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.895 1.86 6.53 1.86 6.53 1.98 6.41 1.98 6.41 1.74 5.35 1.74 5.35 1.42 5.47 1.42 5.47 1.62 6.775 1.62 6.775 0.74 6.51 0.74 6.51 0.5 6.63 0.5 6.63 0.62 6.895 0.62 ;
      POLYGON 5.49 0.74 5.37 0.74 5.37 0.62 4.77 0.62 4.77 1.76 5.11 1.76 5.11 1.8 5.23 1.8 5.23 1.92 4.99 1.92 4.99 1.88 4.65 1.88 4.65 0.62 3.09 0.62 3.09 0.54 2.97 0.54 2.97 0.42 3.21 0.42 3.21 0.5 5.49 0.5 ;
      POLYGON 3.71 1.24 3.59 1.24 3.59 1.12 3.19 1.12 3.19 1.88 2.61 1.88 2.61 1.76 3.07 1.76 3.07 1.12 2.53 1.12 2.53 0.68 2.65 0.68 2.65 1 3.71 1 ;
      POLYGON 2.09 1.4 1.97 1.4 1.97 1.14 1.07 1.14 1.07 1.82 0.95 1.82 0.95 0.68 1.07 0.68 1.07 1.02 2.09 1.02 ;
      POLYGON 1.95 0.54 1.83 0.54 1.83 0.62 1.19 0.62 1.19 0.56 0.78 0.56 0.78 0.68 0.675 0.68 0.675 1.675 0.555 1.675 0.555 0.56 0.66 0.56 0.66 0.44 1.31 0.44 1.31 0.5 1.71 0.5 1.71 0.42 1.95 0.42 ;
  END
END MXI3X2

MACRO AOI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X2 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.11 0.99 4.35 1.11 ;
        RECT 3.205 0.935 4.23 1.055 ;
        RECT 3.005 0.99 3.465 1.09 ;
        RECT 3.005 0.99 3.325 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.42 0.82 2.54 1.15 ;
        RECT 2.39 0.82 2.54 1.145 ;
        RECT 0.525 0.82 2.54 0.94 ;
        RECT 0.525 0.82 0.645 1.15 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.705 1.195 3.99 1.435 ;
        RECT 3.84 1.175 3.99 1.435 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 0.805 1.06 2.22 1.18 ;
        RECT 2.08 1.175 2.25 1.3 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.315 1.3 1.555 1.42 ;
        RECT 1.175 1.52 1.435 1.67 ;
        RECT 1.315 1.3 1.435 1.67 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.965 1.555 4.085 2.01 ;
        RECT 3.125 1.555 4.085 1.675 ;
        RECT 1.54 0.58 3.725 0.7 ;
        RECT 3.125 1.52 3.245 2.01 ;
        RECT 2.625 1.52 3.245 1.64 ;
        RECT 2.625 1.52 2.885 1.67 ;
        RECT 2.765 0.58 2.885 1.67 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 4.185 -0.18 4.305 0.64 ;
        RECT 2.685 0.34 2.925 0.46 ;
        RECT 2.685 -0.18 2.805 0.46 ;
        RECT 0.325 0.46 0.565 0.58 ;
        RECT 0.325 -0.18 0.445 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 2.225 2.03 2.465 2.15 ;
        RECT 2.225 2.03 2.345 2.79 ;
        RECT 1.385 2.03 1.625 2.15 ;
        RECT 1.385 2.03 1.505 2.79 ;
        RECT 0.545 2.03 0.785 2.15 ;
        RECT 0.545 2.03 0.665 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.505 2.25 2.705 2.25 2.705 1.91 1.985 1.91 1.985 2.21 1.865 2.21 1.865 1.91 1.145 1.91 1.145 2.21 1.025 2.21 1.025 1.91 0.305 1.91 0.305 2.21 0.185 2.21 0.185 1.56 0.305 1.56 0.305 1.79 1.865 1.79 1.865 1.56 1.985 1.56 1.985 1.79 2.825 1.79 2.825 2.13 3.545 2.13 3.545 1.795 3.665 1.795 3.665 2.13 4.385 2.13 4.385 1.56 4.505 1.56 ;
  END
END AOI32X2

MACRO OAI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2XL 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.8 0.8 1.145 ;
        RECT 0.61 1 0.73 1.345 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 1.04 1.09 1.525 ;
        RECT 0.94 1.04 1.09 1.495 ;
    END
  END A0N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.13 2.83 1.6 ;
        RECT 2.68 1.1 2.8 1.6 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.11 3.41 1.435 ;
        RECT 3.19 1.28 3.31 1.6 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.192 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.95 0.89 3.07 1.84 ;
        RECT 2.92 0.68 3.04 1.01 ;
        RECT 2.625 1.72 3.07 1.84 ;
        RECT 2.44 1.84 2.885 1.96 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 1.96 -0.18 2.08 0.92 ;
        RECT 0.61 -0.18 0.73 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.08 1.96 3.32 2.08 ;
        RECT 3.08 1.96 3.2 2.79 ;
        RECT 1.86 1.9 1.98 2.79 ;
        RECT 0.79 1.645 0.91 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.46 0.92 3.34 0.92 3.34 0.56 2.68 0.56 2.68 0.8 2.62 0.8 2.62 0.92 2.56 0.92 2.56 1.4 1.48 1.4 1.48 0.68 1.6 0.68 1.6 1.28 2.44 1.28 2.44 0.8 2.5 0.8 2.5 0.68 2.56 0.68 2.56 0.44 3.46 0.44 ;
      POLYGON 2.44 0.52 2.32 0.52 2.32 1.16 1.72 1.16 1.72 0.56 0.97 0.56 0.97 0.68 0.255 0.68 0.255 1.525 0.49 1.525 0.49 1.765 0.37 1.765 0.37 1.645 0.135 1.645 0.135 0.56 0.85 0.56 0.85 0.44 1.84 0.44 1.84 1.04 2.2 1.04 2.2 0.4 2.44 0.4 ;
      POLYGON 1.86 1.64 1.33 1.64 1.33 1.765 1.21 1.765 1.21 0.92 1.09 0.92 1.09 0.68 1.21 0.68 1.21 0.8 1.33 0.8 1.33 1.52 1.86 1.52 ;
  END
END OAI2BB2XL

MACRO SMDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX1 0 0 ;
  SIZE 10.15 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.22 0.895 1.46 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.34 0.8 1.725 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.095 1.2 6.215 1.44 ;
        RECT 5.87 1.2 6.215 1.435 ;
        RECT 5.87 1.175 6.02 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.595 0.995 7.76 1.435 ;
        RECT 7.595 0.975 7.715 1.44 ;
    END
  END SE
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.9 1 8.055 1.45 ;
        RECT 7.935 0.975 8.055 1.45 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.21 9.555 1.465 ;
        RECT 9.255 1.22 9.555 1.45 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.675 0.97 9.795 1.21 ;
        RECT 8.645 0.97 9.795 1.09 ;
        RECT 9.005 0.94 9.265 1.09 ;
        RECT 8.915 0.97 9.155 1.1 ;
        RECT 8.415 1.01 8.765 1.13 ;
        RECT 8.415 1.01 8.535 1.44 ;
    END
  END S0
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.15 0.18 ;
        RECT 9.475 -0.18 9.595 0.82 ;
        RECT 8.165 -0.18 8.285 0.65 ;
        RECT 6.175 -0.18 6.295 0.8 ;
        RECT 3.905 -0.18 4.145 0.36 ;
        RECT 1.785 0.5 2.025 0.62 ;
        RECT 1.785 -0.18 1.905 0.62 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.15 2.79 ;
        RECT 9.385 1.825 9.505 2.79 ;
        RECT 7.935 1.85 8.055 2.79 ;
        RECT 6.085 1.85 6.205 2.79 ;
        RECT 3.905 2 4.145 2.12 ;
        RECT 3.905 2 4.025 2.79 ;
        RECT 1.925 2 2.165 2.12 ;
        RECT 1.925 2 2.045 2.79 ;
        RECT 0.555 1.845 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.035 1.705 9.985 1.705 9.985 1.825 9.865 1.825 9.865 1.705 8.885 1.705 8.885 1.24 9.005 1.24 9.005 1.585 9.915 1.585 9.915 0.85 9.895 0.85 9.895 0.58 10.015 0.58 10.015 0.73 10.035 0.73 ;
      POLYGON 8.955 0.83 8.525 0.83 8.525 0.89 8.295 0.89 8.295 1.57 8.575 1.57 8.575 1.56 8.695 1.56 8.695 2.21 8.575 2.21 8.575 1.69 7.325 1.69 7.325 1.82 7.205 1.82 7.205 1.56 7.355 1.56 7.355 0.84 7.295 0.84 7.295 0.6 7.415 0.6 7.415 0.72 7.475 0.72 7.475 1.57 8.175 1.57 8.175 0.77 8.405 0.77 8.405 0.71 8.835 0.71 8.835 0.58 8.955 0.58 ;
      POLYGON 7.805 0.84 7.685 0.84 7.685 0.6 7.585 0.6 7.585 0.48 7.175 0.48 7.175 0.96 7.235 0.96 7.235 1.44 7.085 1.44 7.085 1.97 7.635 1.97 7.635 2.21 7.515 2.21 7.515 2.09 6.965 2.09 6.965 1.44 6.575 1.44 6.575 1.2 6.695 1.2 6.695 1.32 7.115 1.32 7.115 1.08 7.055 1.08 7.055 0.36 7.705 0.36 7.705 0.48 7.805 0.48 ;
      POLYGON 6.935 1.04 6.455 1.04 6.455 1.56 6.845 1.56 6.845 2.21 6.725 2.21 6.725 1.68 5.425 1.68 5.425 1.64 5.305 1.64 5.305 1.52 5.425 1.52 5.425 0.72 5.305 0.72 5.305 0.6 5.545 0.6 5.545 1.56 6.335 1.56 6.335 0.92 6.815 0.92 6.815 0.62 6.935 0.62 ;
      POLYGON 5.875 0.8 5.755 0.8 5.755 0.48 5.185 0.48 5.185 1.12 5.205 1.12 5.205 1.36 5.185 1.36 5.185 1.8 5.725 1.8 5.725 1.91 5.845 1.91 5.845 2.03 5.605 2.03 5.605 1.92 5.065 1.92 5.065 0.48 4.585 0.48 4.585 0.92 4.705 0.92 4.705 1.04 4.465 1.04 4.465 0.6 3.665 0.6 3.665 0.48 3.185 0.48 3.185 0.96 3.405 0.96 3.405 1.2 3.285 1.2 3.285 1.08 3.065 1.08 3.065 0.36 3.785 0.36 3.785 0.48 4.465 0.48 4.465 0.36 5.875 0.36 ;
      POLYGON 4.945 1.98 4.825 1.98 4.825 1.28 3.765 1.28 3.765 1.16 4.825 1.16 4.825 0.72 4.705 0.72 4.705 0.6 4.945 0.6 ;
      POLYGON 4.725 2.24 4.37 2.24 4.37 1.88 3.165 1.88 3.165 2.22 2.36 2.22 2.36 1.88 1.035 1.88 1.035 0.68 1.155 0.68 1.155 1.76 2.36 1.76 2.36 1.1 2.285 1.1 2.285 0.98 2.525 0.98 2.525 1.1 2.48 1.1 2.48 2.1 3.045 2.1 3.045 1.32 2.885 1.32 2.885 1.2 3.165 1.2 3.165 1.76 4.49 1.76 4.49 2.12 4.725 2.12 ;
      POLYGON 4.345 1.04 3.645 1.04 3.645 1.64 3.405 1.64 3.405 1.52 3.525 1.52 3.525 0.84 3.305 0.84 3.305 0.6 3.545 0.6 3.545 0.72 3.645 0.72 3.645 0.92 4.345 0.92 ;
      POLYGON 2.925 1.98 2.805 1.98 2.805 1.56 2.645 1.56 2.645 0.78 2.265 0.78 2.265 0.86 1.785 0.86 1.785 1.12 1.665 1.12 1.665 0.74 2.145 0.74 2.145 0.66 2.645 0.66 2.645 0.54 2.765 0.54 2.765 1.44 2.925 1.44 ;
      POLYGON 2.165 1.3 2.025 1.3 2.025 1.36 1.545 1.36 1.545 1.52 1.685 1.52 1.685 1.64 1.425 1.64 1.425 0.56 0.915 0.56 0.915 1.1 0.535 1.1 0.535 1.24 0.415 1.24 0.415 0.98 0.795 0.98 0.795 0.44 1.545 0.44 1.545 1.24 1.905 1.24 1.905 1.18 2.165 1.18 ;
  END
END SMDFFHQX1

MACRO MXI4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.6133 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 1.2 1.155 1.44 ;
        RECT 0.39 1.2 1.155 1.32 ;
        RECT 0.36 1.465 0.51 1.725 ;
        RECT 0.39 1.2 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.44 0.835 1.85 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.115 1.29 2.255 1.685 ;
        RECT 2.08 1.34 2.25 1.725 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.31 2.615 1.725 ;
        RECT 2.495 1.29 2.615 1.725 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 1.36 4.005 1.725 ;
        RECT 3.835 1.28 3.97 1.65 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6952 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.715 1.57 7.955 1.69 ;
        RECT 6.755 0.95 7.955 1.07 ;
        RECT 7.835 0.6 7.955 1.07 ;
        RECT 7.715 0.95 7.835 1.69 ;
        RECT 7.61 0.95 7.835 1.435 ;
        RECT 6.755 1.57 6.995 1.69 ;
        RECT 6.855 0.95 6.975 1.69 ;
        RECT 6.755 0.6 6.875 1.07 ;
    END
  END Y
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.135 1.52 8.655 1.64 ;
        RECT 7.48 1.81 8.395 1.93 ;
        RECT 8.275 1.52 8.395 1.93 ;
        RECT 8.135 1.52 8.395 1.67 ;
        RECT 7.48 1.81 7.6 2.17 ;
        RECT 5.89 2.05 7.6 2.17 ;
        RECT 4.575 2.13 6.01 2.25 ;
        RECT 4.575 1.33 4.695 2.25 ;
    END
  END S1
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.315 -0.18 8.435 0.84 ;
        RECT 7.235 0.47 7.475 0.59 ;
        RECT 7.355 -0.18 7.475 0.59 ;
        RECT 6.275 -0.18 6.395 0.79 ;
        RECT 4.085 -0.18 4.205 0.92 ;
        RECT 2.355 -0.18 2.475 0.38 ;
        RECT 0.495 0.72 0.735 0.84 ;
        RECT 0.495 -0.18 0.615 0.84 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.195 2.05 8.435 2.17 ;
        RECT 8.195 2.05 8.315 2.79 ;
        RECT 7.235 2.29 7.475 2.79 ;
        RECT 6.13 2.29 6.37 2.79 ;
        RECT 3.7 2.085 3.94 2.205 ;
        RECT 3.7 2.085 3.82 2.79 ;
        RECT 2.055 2.085 2.295 2.205 ;
        RECT 2.055 2.085 2.175 2.79 ;
        RECT 0.715 1.97 0.835 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.895 1.88 8.855 1.88 8.855 2.04 8.735 2.04 8.735 1.76 8.775 1.76 8.775 1.08 8.075 1.08 8.075 0.48 7.715 0.48 7.715 0.83 6.995 0.83 6.995 0.48 6.635 0.48 6.635 1.69 5.435 1.69 5.435 1.54 4.895 1.54 4.895 1.02 5.015 1.02 5.015 1.42 5.435 1.42 5.435 1.3 5.555 1.3 5.555 1.57 6.515 1.57 6.515 0.36 7.115 0.36 7.115 0.71 7.595 0.71 7.595 0.36 8.195 0.36 8.195 0.96 8.605 0.96 8.605 0.72 8.735 0.72 8.735 0.6 8.855 0.6 8.855 0.72 8.895 0.72 ;
      POLYGON 7.235 1.93 5.315 1.93 5.315 2.01 5.195 2.01 5.195 1.67 5.315 1.67 5.315 1.81 7.115 1.81 7.115 1.43 7.095 1.43 7.095 1.19 7.215 1.19 7.215 1.31 7.235 1.31 ;
      POLYGON 6.395 1.45 5.675 1.45 5.675 1.01 5.135 1.01 5.135 0.89 4.955 0.89 4.955 0.65 5.075 0.65 5.075 0.77 5.255 0.77 5.255 0.89 5.795 0.89 5.795 1.33 6.275 1.33 6.275 1.19 6.395 1.19 ;
      POLYGON 6.035 1.21 5.915 1.21 5.915 0.53 4.445 0.53 4.445 1.16 3.715 1.16 3.715 1.725 3.34 1.725 3.34 2.01 2.915 2.01 2.915 1.89 3.22 1.89 3.22 1.605 3.595 1.605 3.595 0.9 3.255 0.9 3.255 0.86 3.135 0.86 3.135 0.74 3.375 0.74 3.375 0.78 3.715 0.78 3.715 1.04 4.325 1.04 4.325 0.41 6.035 0.41 ;
      POLYGON 4.375 1.965 3.58 1.965 3.58 2.25 2.665 2.25 2.665 1.97 2.415 1.97 2.415 1.965 1.74 1.965 1.74 1.97 1.475 1.97 1.475 2.09 1.355 2.09 1.355 1.97 1.275 1.97 1.275 0.66 1.395 0.66 1.395 1.85 1.62 1.85 1.62 1.845 2.535 1.845 2.535 1.85 2.785 1.85 2.785 2.13 3.46 2.13 3.46 1.845 4.255 1.845 4.255 1.33 4.375 1.33 ;
      POLYGON 3.475 1.26 3.355 1.26 3.355 1.17 2.935 1.17 2.935 1.73 2.815 1.73 2.815 1.17 1.995 1.17 1.995 1.18 1.755 1.18 1.755 1.05 3.355 1.05 3.355 1.02 3.475 1.02 ;
      POLYGON 3.035 0.62 1.635 0.62 1.635 1.725 1.515 1.725 1.515 0.54 0.975 0.54 0.975 1.08 0.24 1.08 0.24 1.85 0.355 1.85 0.355 2.09 0.235 2.09 0.235 1.97 0.12 1.97 0.12 0.78 0.135 0.78 0.135 0.66 0.255 0.66 0.255 0.96 0.855 0.96 0.855 0.42 0.995 0.42 0.995 0.4 1.235 0.4 1.235 0.42 1.635 0.42 1.635 0.5 2.915 0.5 2.915 0.36 3.035 0.36 ;
  END
END MXI4X4

MACRO DFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQXL 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 1.465 0.855 1.725 ;
        RECT 0.665 1.385 0.855 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.965 1.49 5.27 1.665 ;
        RECT 4.89 1.52 5.205 1.72 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.965 ;
        RECT 0.07 1.465 0.255 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.025 0.67 5.265 0.79 ;
        RECT 5.025 -0.18 5.145 0.79 ;
        RECT 3.605 0.43 3.845 0.55 ;
        RECT 3.605 -0.18 3.725 0.55 ;
        RECT 1.905 -0.18 2.025 0.86 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.105 1.87 5.225 2.79 ;
        RECT 3.505 2.29 3.745 2.79 ;
        RECT 1.785 2.29 2.025 2.79 ;
        RECT 0.555 1.845 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.685 1.51 5.645 1.51 5.645 1.99 5.525 1.99 5.525 1.39 5.565 1.39 5.565 1.03 4.785 1.03 4.785 0.5 4.085 0.5 4.085 0.79 3.365 0.79 3.365 0.5 3.005 0.5 3.005 1.15 3.205 1.15 3.205 1.27 2.665 1.27 2.665 1.53 2.585 1.53 2.585 1.65 2.465 1.65 2.465 1.41 2.545 1.41 2.545 1.15 2.885 1.15 2.885 0.38 3.485 0.38 3.485 0.67 3.965 0.67 3.965 0.38 4.165 0.38 4.165 0.36 4.405 0.36 4.405 0.38 4.905 0.38 4.905 0.91 5.565 0.91 5.565 0.62 5.685 0.62 ;
      POLYGON 5.445 1.27 5.325 1.27 5.325 1.37 4.785 1.37 4.785 1.4 4.685 1.4 4.685 2.17 2.905 2.17 2.905 2.25 2.145 2.25 2.145 2.17 0.975 2.17 0.975 1.725 1.035 1.725 1.035 0.68 1.155 0.68 1.155 1.845 1.095 1.845 1.095 2.05 2.265 2.05 2.265 2.13 2.785 2.13 2.785 1.55 2.825 1.55 2.825 1.43 2.945 1.43 2.945 1.67 2.905 1.67 2.905 2.05 4.565 2.05 4.565 1.65 4.105 1.65 4.105 1.41 4.225 1.41 4.225 1.53 4.565 1.53 4.565 1.25 4.665 1.25 4.665 1.16 4.785 1.16 4.785 1.25 5.205 1.25 5.205 1.15 5.445 1.15 ;
      POLYGON 4.505 0.86 4.325 0.86 4.325 1.29 3.985 1.29 3.985 1.77 4.325 1.77 4.325 1.81 4.445 1.81 4.445 1.93 4.205 1.93 4.205 1.89 3.865 1.89 3.865 1.5 3.685 1.5 3.685 1.62 3.565 1.62 3.565 1.38 3.865 1.38 3.865 1.17 4.205 1.17 4.205 0.74 4.385 0.74 4.385 0.62 4.505 0.62 ;
      POLYGON 3.745 1.26 3.445 1.26 3.445 1.93 3.025 1.93 3.025 1.81 3.325 1.81 3.325 1.03 3.125 1.03 3.125 0.62 3.245 0.62 3.245 0.91 3.445 0.91 3.445 1.14 3.625 1.14 3.625 1.02 3.745 1.02 ;
      POLYGON 2.765 0.8 2.345 0.8 2.345 1.77 2.665 1.77 2.665 2.01 2.545 2.01 2.545 1.89 2.225 1.89 2.225 1.65 1.745 1.65 1.745 1.41 1.865 1.41 1.865 1.53 2.225 1.53 2.225 0.68 2.765 0.68 ;
      POLYGON 2.105 1.31 1.985 1.31 1.985 1.29 1.605 1.29 1.605 1.93 1.305 1.93 1.305 1.81 1.485 1.81 1.485 0.56 0.915 0.56 0.915 1.16 0.515 1.16 0.515 1.28 0.395 1.28 0.395 1.04 0.795 1.04 0.795 0.44 1.605 0.44 1.605 1.17 1.985 1.17 1.985 1.07 2.105 1.07 ;
  END
END DFFQXL

MACRO TLATSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX2 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.01 3.7 1.48 ;
        RECT 3.565 0.98 3.685 1.48 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.16 0.835 1.58 ;
        RECT 0.65 1.16 0.835 1.565 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.33 3.12 1.725 ;
        RECT 2.88 1.33 3.12 1.45 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.625 1.215 4.915 1.43 ;
        RECT 4.625 1.095 4.745 1.47 ;
    END
  END SN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.525 0.94 5.785 1.09 ;
        RECT 5.285 0.94 5.785 1.06 ;
        RECT 5.285 0.615 5.405 1.335 ;
        RECT 5.185 1.215 5.305 2.11 ;
        RECT 5.185 0.495 5.305 0.735 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.885 0.885 7.18 1.145 ;
        RECT 6.885 0.765 7.005 1.58 ;
        RECT 6.865 1.46 6.985 2.11 ;
        RECT 6.865 0.595 6.985 0.885 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 7.285 -0.18 7.405 0.645 ;
        RECT 6.445 -0.18 6.565 0.645 ;
        RECT 5.605 -0.18 5.725 0.645 ;
        RECT 4.765 -0.18 4.885 0.735 ;
        RECT 2.715 0.61 2.955 0.73 ;
        RECT 2.835 -0.18 2.955 0.73 ;
        RECT 0.495 0.68 0.735 0.8 ;
        RECT 0.495 -0.18 0.615 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 7.285 1.46 7.405 2.79 ;
        RECT 6.445 1.46 6.565 2.79 ;
        RECT 5.605 1.46 5.725 2.79 ;
        RECT 4.765 1.59 4.885 2.79 ;
        RECT 3.865 2.23 3.985 2.79 ;
        RECT 3.145 2.23 3.265 2.79 ;
        RECT 2.245 2.29 2.485 2.79 ;
        RECT 0.715 1.94 0.835 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.765 1.24 6.145 1.24 6.145 2.11 6.025 2.11 6.025 0.595 6.145 0.595 6.145 1.12 6.765 1.12 ;
      POLYGON 5.165 1.095 4.925 1.095 4.925 0.975 4.465 0.975 4.465 2.11 4.345 2.11 4.345 0.975 4.125 0.975 4.125 0.5 3.195 0.5 3.195 0.97 2.275 0.97 2.275 0.48 2.155 0.48 2.155 0.36 2.395 0.36 2.395 0.85 3.075 0.85 3.075 0.38 4.245 0.38 4.245 0.855 5.165 0.855 ;
      POLYGON 4.185 2.11 2.41 2.11 2.41 2.17 1.495 2.17 1.495 1.75 1.615 1.75 1.615 1.57 1.655 1.57 1.655 0.62 1.775 0.62 1.775 1.69 1.735 1.69 1.735 1.87 1.615 1.87 1.615 2.05 2.29 2.05 2.29 1.99 4.065 1.99 4.065 1.27 4.185 1.27 ;
      POLYGON 3.94 1.72 3.625 1.72 3.625 1.84 3.505 1.84 3.505 1.72 3.24 1.72 3.24 1.21 1.915 1.21 1.915 0.5 1.535 0.5 1.535 1.45 1.415 1.45 1.415 1.04 0.515 1.04 0.515 1.2 0.395 1.2 0.395 0.92 1.415 0.92 1.415 0.38 2.035 0.38 2.035 0.96 2.095 0.96 2.095 1.09 3.36 1.09 3.36 1.6 3.82 1.6 3.82 0.86 3.475 0.86 3.475 0.62 3.595 0.62 3.595 0.74 3.94 0.74 ;
      POLYGON 2.845 1.87 2.095 1.87 2.095 1.93 1.855 1.93 1.855 1.81 1.975 1.81 1.975 1.75 2.845 1.75 ;
      POLYGON 1.235 1.28 1.075 1.28 1.075 1.82 0.355 1.82 0.355 1.99 0.235 1.99 0.235 1.87 0.155 1.87 0.155 0.86 0.135 0.86 0.135 0.62 0.255 0.62 0.255 0.74 0.275 0.74 0.275 1.7 0.955 1.7 0.955 1.16 1.235 1.16 ;
  END
END TLATSRX2

MACRO SDFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX2 0 0 ;
  SIZE 13.34 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.08 1.045 2.32 1.25 ;
        RECT 2.1 1.045 2.25 1.435 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.27 2.13 7.47 2.25 ;
        RECT 6.27 1.7 6.39 2.25 ;
        RECT 5.67 1.7 6.39 1.82 ;
        RECT 4.59 2.13 5.79 2.25 ;
        RECT 5.67 1.7 5.79 2.25 ;
        RECT 4.35 2.08 4.71 2.2 ;
        RECT 4.35 1.4 4.47 2.2 ;
        RECT 2.88 1.4 4.47 1.52 ;
        RECT 2.88 1.23 3 1.52 ;
        RECT 2.68 1.195 2.92 1.38 ;
        RECT 2.625 1.23 3 1.38 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.535 1.16 10.655 1.4 ;
        RECT 10.165 1.23 10.655 1.38 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.895 0.94 11.015 1.305 ;
        RECT 10.8 0.785 10.95 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 1.23 12.455 1.43 ;
        RECT 12.075 1.245 12.455 1.42 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.83 1.175 12.98 1.435 ;
        RECT 12.695 0.99 12.95 1.23 ;
        RECT 11.375 0.99 12.95 1.11 ;
        RECT 11.875 0.98 12.115 1.11 ;
        RECT 11.375 0.99 11.495 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 1.755 0.8 2.015 ;
        RECT 0.63 1.54 0.77 2.015 ;
        RECT 0.63 1.54 0.75 2.19 ;
        RECT 0.59 0.8 0.71 1.66 ;
        RECT 0.57 0.68 0.69 0.92 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.34 0.18 ;
        RECT 12.435 -0.18 12.555 0.84 ;
        RECT 10.915 -0.18 11.155 0.32 ;
        RECT 9.94 -0.18 10.18 0.32 ;
        RECT 7.79 -0.18 7.91 0.64 ;
        RECT 2.4 -0.18 2.52 0.685 ;
        RECT 0.99 -0.18 1.11 0.74 ;
        RECT 0.15 -0.18 0.27 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.34 2.79 ;
        RECT 12.215 1.795 12.335 2.79 ;
        RECT 10.895 1.56 11.015 2.79 ;
        RECT 10 1.76 10.12 2.79 ;
        RECT 7.63 1.88 7.87 2 ;
        RECT 7.63 1.88 7.75 2.79 ;
        RECT 6.03 1.94 6.15 2.79 ;
        RECT 5.91 1.94 6.15 2.06 ;
        RECT 3.66 1.88 3.9 2 ;
        RECT 3.68 1.88 3.8 2.79 ;
        RECT 2.4 1.795 2.52 2.79 ;
        RECT 2.28 1.795 2.52 1.915 ;
        RECT 1.05 1.54 1.17 2.79 ;
        RECT 0.21 1.54 0.33 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.22 1.975 12.575 1.975 12.575 1.855 13.1 1.855 13.1 1.675 11.835 1.675 11.835 1.42 11.655 1.42 11.655 1.3 11.955 1.3 11.955 1.555 13.1 1.555 13.1 0.87 12.855 0.87 12.855 0.6 12.975 0.6 12.975 0.75 13.22 0.75 ;
      POLYGON 11.855 0.665 11.255 0.665 11.255 1.56 11.655 1.56 11.655 2.21 11.535 2.21 11.535 1.68 11.135 1.68 11.135 0.665 10.87 0.665 10.87 0.56 8.97 0.56 8.97 0.9 9.21 0.9 9.21 1.54 9.31 1.54 9.31 1.77 9.07 1.77 9.07 1.54 9.09 1.54 9.09 1.02 8.85 1.02 8.85 0.44 10.99 0.44 10.99 0.545 11.855 0.545 ;
      POLYGON 10.655 1.74 10.415 1.74 10.415 1.64 9.88 1.64 9.88 2.25 7.99 2.25 7.99 1.76 7.51 1.76 7.51 2.01 6.51 2.01 6.51 1.58 5.55 1.58 5.55 2.01 4.83 2.01 4.83 1.26 4.85 1.26 4.85 0.84 4.95 0.84 4.95 0.48 4.47 0.48 4.47 1.04 4.23 1.04 4.23 0.92 4.35 0.92 4.35 0.36 5.07 0.36 5.07 0.96 4.97 0.96 4.97 1.38 4.95 1.38 4.95 1.89 5.43 1.89 5.43 1.46 6.63 1.46 6.63 1.89 7.39 1.89 7.39 1.64 8.11 1.64 8.11 2.13 9.76 2.13 9.76 1.52 9.8 1.52 9.8 0.92 10.335 0.92 10.335 0.68 10.575 0.68 10.575 0.8 10.455 0.8 10.455 1.04 9.92 1.04 9.92 1.52 10.535 1.52 10.535 1.62 10.655 1.62 ;
      POLYGON 9.7 0.8 9.64 0.8 9.64 2.01 8.23 2.01 8.23 1.16 7.75 1.16 7.75 1.28 6.99 1.28 6.99 1.1 5.55 1.1 5.55 1.04 5.43 1.04 5.43 0.92 5.67 0.92 5.67 0.98 7.11 0.98 7.11 1.16 7.63 1.16 7.63 1.04 8.23 1.04 8.23 1 8.47 1 8.47 1.12 8.35 1.12 8.35 1.89 8.83 1.89 8.83 1.14 8.97 1.14 8.97 1.38 8.95 1.38 8.95 1.89 9.52 1.89 9.52 0.8 9.46 0.8 9.46 0.68 9.7 0.68 ;
      POLYGON 8.71 1.77 8.47 1.77 8.47 1.6 8.59 1.6 8.59 0.74 8.285 0.74 8.285 0.88 7.755 0.88 7.755 0.92 7.47 0.92 7.47 1.04 7.23 1.04 7.23 0.92 7.35 0.92 7.35 0.8 7.635 0.8 7.635 0.76 8.165 0.76 8.165 0.62 8.43 0.62 8.43 0.5 8.55 0.5 8.55 0.62 8.71 0.62 ;
      POLYGON 8.11 1.4 7.99 1.4 7.99 1.52 7.27 1.52 7.27 1.77 7.15 1.77 7.15 1.52 6.75 1.52 6.75 1.34 5.31 1.34 5.31 1.77 5.07 1.77 5.07 1.5 5.19 1.5 5.19 0.54 5.31 0.54 5.31 0.68 6.155 0.68 6.155 0.74 6.83 0.74 6.83 0.6 7.13 0.6 7.13 0.72 6.95 0.72 6.95 0.86 6.035 0.86 6.035 0.8 5.31 0.8 5.31 1.22 6.87 1.22 6.87 1.4 7.87 1.4 7.87 1.28 8.11 1.28 ;
      POLYGON 7.49 0.68 7.37 0.68 7.37 0.48 6.71 0.48 6.71 0.62 6.47 0.62 6.47 0.5 6.59 0.5 6.59 0.36 7.49 0.36 ;
      POLYGON 4.83 0.72 4.71 0.72 4.71 1.96 4.59 1.96 4.59 1.28 3.12 1.28 3.12 1.075 2.69 1.075 2.69 0.925 2.16 0.925 2.16 0.48 1.35 0.48 1.35 1.18 1.23 1.18 1.23 0.36 2.28 0.36 2.28 0.805 2.81 0.805 2.81 0.955 3.24 0.955 3.24 1.16 4.59 1.16 4.59 0.6 4.83 0.6 ;
      POLYGON 4.23 0.72 4.11 0.72 4.11 0.925 3.36 0.925 3.36 0.725 3.18 0.725 3.18 0.605 3.48 0.605 3.48 0.805 3.99 0.805 3.99 0.6 4.23 0.6 ;
      POLYGON 4.23 1.96 4.11 1.96 4.11 1.76 3 1.76 3 1.975 2.88 1.975 2.88 1.64 4.23 1.64 ;
      POLYGON 3.78 0.685 3.66 0.685 3.66 0.485 2.94 0.485 2.94 0.685 2.82 0.685 2.82 0.365 3.78 0.365 ;
      POLYGON 3.56 2.25 3.055 2.25 3.055 2.215 2.64 2.215 2.64 1.675 1.86 1.675 1.86 1.55 1.84 1.55 1.84 0.72 1.8 0.72 1.8 0.6 2.04 0.6 2.04 0.72 1.96 0.72 1.96 1.43 1.98 1.43 1.98 1.555 2.76 1.555 2.76 2.095 3.175 2.095 3.175 2.13 3.56 2.13 ;
      POLYGON 2.28 2.25 2.04 2.25 2.04 2.18 1.47 2.18 1.47 1.42 0.83 1.42 0.83 1.18 0.95 1.18 0.95 1.3 1.47 1.3 1.47 0.6 1.59 0.6 1.59 2.06 2.16 2.06 2.16 2.13 2.28 2.13 ;
  END
END SDFFSRHQX2

MACRO SEDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX1 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.33 0.76 1.45 1.15 ;
        RECT 0.59 0.76 1.45 0.88 ;
        RECT 0.445 1.07 0.71 1.19 ;
        RECT 0.59 0.76 0.71 1.19 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.445 1.07 0.565 1.38 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.91 1.02 1.09 1.44 ;
        RECT 0.91 1 1.03 1.44 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.165 ;
        RECT 2.71 0.94 2.83 1.34 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 1.225 4.625 1.46 ;
        RECT 4.32 1.13 4.56 1.345 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.8 1.03 10.95 1.5 ;
        RECT 10.8 1.03 10.92 1.53 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.9 0.68 6.02 1.025 ;
        RECT 5.895 0.905 6.015 1.99 ;
        RECT 5.58 1.025 6.015 1.145 ;
        RECT 5.58 0.885 5.73 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.615 -0.18 10.735 0.67 ;
        RECT 8.625 0.43 8.865 0.55 ;
        RECT 8.625 -0.18 8.745 0.55 ;
        RECT 6.905 0.41 7.145 0.53 ;
        RECT 6.905 -0.18 7.025 0.53 ;
        RECT 5.36 -0.18 5.6 0.32 ;
        RECT 4.46 -0.18 4.58 0.64 ;
        RECT 2.31 0.46 2.55 0.58 ;
        RECT 2.31 -0.18 2.43 0.58 ;
        RECT 0.83 -0.18 0.95 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.635 1.89 10.755 2.79 ;
        RECT 8.405 2.25 8.645 2.79 ;
        RECT 6.805 1.49 6.925 2.79 ;
        RECT 5.475 1.34 5.595 2.79 ;
        RECT 4.54 1.9 4.66 2.79 ;
        RECT 2.21 1.7 2.33 2.79 ;
        RECT 0.77 1.8 0.89 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.235 1.95 10.995 1.95 10.995 1.77 10.515 1.77 10.515 2.25 8.965 2.25 8.965 2.13 8.025 2.13 8.025 2.25 7.665 2.25 7.665 2.13 7.905 2.13 7.905 2.01 9.085 2.01 9.085 2.13 10.395 2.13 10.395 1.65 10.56 1.65 10.56 1.03 10.455 1.03 10.455 0.79 10.855 0.79 10.855 0.67 11.035 0.67 11.035 0.43 11.155 0.43 11.155 0.79 10.975 0.79 10.975 0.91 10.68 0.91 10.68 1.65 11.115 1.65 11.115 1.83 11.235 1.83 ;
      POLYGON 10.315 0.67 10.275 0.67 10.275 2.01 9.465 2.01 9.465 1.89 7.685 1.89 7.685 1.25 7.465 1.25 7.465 1.37 7.345 1.37 7.345 1.13 7.905 1.13 7.905 0.86 8.025 0.86 8.025 1.25 7.805 1.25 7.805 1.77 9.465 1.77 9.465 1.33 9.345 1.33 9.345 1.21 9.585 1.21 9.585 1.89 10.155 1.89 10.155 0.55 10.195 0.55 10.195 0.43 10.315 0.43 ;
      POLYGON 9.945 1.77 9.705 1.77 9.705 1.53 9.805 1.53 9.805 0.48 9.13 0.48 9.13 0.79 8.385 0.79 8.385 0.48 7.385 0.48 7.385 0.77 6.665 0.77 6.665 0.48 6.145 0.48 6.145 0.56 4.82 0.56 4.82 0.88 4.085 0.88 4.085 0.83 3.94 0.83 3.94 1.77 3.82 1.77 3.82 0.59 3.94 0.59 3.94 0.71 4.205 0.71 4.205 0.76 4.7 0.76 4.7 0.44 6.025 0.44 6.025 0.36 6.785 0.36 6.785 0.65 7.265 0.65 7.265 0.36 8.505 0.36 8.505 0.67 9.01 0.67 9.01 0.36 9.925 0.36 9.925 1.53 9.945 1.53 ;
      POLYGON 9.565 0.72 9.445 0.72 9.445 1.09 9.225 1.09 9.225 1.53 9.345 1.53 9.345 1.65 9.105 1.65 9.105 1.39 8.385 1.39 8.385 1.15 8.505 1.15 8.505 1.27 9.105 1.27 9.105 0.97 9.325 0.97 9.325 0.6 9.565 0.6 ;
      POLYGON 8.845 1.15 8.725 1.15 8.725 1.03 8.265 1.03 8.265 1.65 7.925 1.65 7.925 1.53 8.145 1.53 8.145 0.72 8.025 0.72 8.025 0.6 8.265 0.6 8.265 0.91 8.845 0.91 ;
      POLYGON 7.845 0.72 7.725 0.72 7.725 1.01 7.225 1.01 7.225 1.49 7.565 1.49 7.565 1.99 7.445 1.99 7.445 1.61 7.105 1.61 7.105 1.37 6.525 1.37 6.525 1.13 6.645 1.13 6.645 1.25 7.105 1.25 7.105 0.89 7.605 0.89 7.605 0.6 7.845 0.6 ;
      POLYGON 6.985 1.13 6.865 1.13 6.865 1.01 6.405 1.01 6.405 1.99 6.285 1.99 6.285 1.24 6.14 1.24 6.14 0.89 6.285 0.89 6.285 0.6 6.545 0.6 6.545 0.72 6.405 0.72 6.405 0.89 6.985 0.89 ;
      POLYGON 5.175 1.78 4.42 1.78 4.42 2.25 2.45 2.25 2.45 1.58 2.19 1.58 2.19 1.24 2.31 1.24 2.31 1.46 2.57 1.46 2.57 2.13 4.3 2.13 4.3 1.66 5.055 1.66 5.055 1.22 4.94 1.22 4.94 0.68 5.06 0.68 5.06 1.1 5.175 1.1 ;
      POLYGON 4.18 2.01 2.69 2.01 2.69 1.46 3.005 1.46 3.005 0.77 2.91 0.77 2.91 0.65 3.15 0.65 3.15 0.77 3.125 0.77 3.125 1.58 2.81 1.58 2.81 1.89 3.58 1.89 3.58 1.17 3.52 1.17 3.52 0.93 3.7 0.93 3.7 1.89 4.06 1.89 4.06 1.15 4.18 1.15 ;
      POLYGON 3.48 0.77 3.4 0.77 3.4 1.49 3.46 1.49 3.46 1.77 3.34 1.77 3.34 1.61 3.28 1.61 3.28 0.65 3.36 0.65 3.36 0.53 2.79 0.53 2.79 0.82 1.73 0.82 1.73 0.83 1.69 0.83 1.69 2.01 1.57 2.01 1.57 0.71 1.61 0.71 1.61 0.59 1.73 0.59 1.73 0.7 2.67 0.7 2.67 0.41 3.48 0.41 ;
      POLYGON 2.05 1.09 1.93 1.09 1.93 2.25 1.33 2.25 1.33 1.8 1.21 1.8 1.21 1.68 0.41 1.68 0.41 1.8 0.29 1.8 0.29 1.68 0.065 1.68 0.065 0.83 0.35 0.83 0.35 0.59 0.47 0.59 0.47 0.95 0.185 0.95 0.185 1.56 1.21 1.56 1.21 1.3 1.45 1.3 1.45 1.42 1.33 1.42 1.33 1.68 1.45 1.68 1.45 2.13 1.81 2.13 1.81 0.97 2.05 0.97 ;
  END
END SEDFFHQX1

MACRO MX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.58 1.155 1.7 ;
        RECT 1.035 1.12 1.155 1.7 ;
        RECT 0.36 1.465 0.51 1.725 ;
        RECT 0.375 1.46 0.495 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.02 0.815 1.46 ;
        RECT 0.695 1 0.815 1.46 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.21 2.015 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 1.175 2.54 1.435 ;
        RECT 2.315 1.055 2.435 2.21 ;
        RECT 2.255 0.59 2.375 1.175 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.835 -0.18 1.955 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.895 1.6 2.015 2.79 ;
        RECT 0.555 1.92 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.135 1.09 1.635 1.09 1.635 1.94 1.375 1.94 1.375 1.98 1.135 1.98 1.135 1.86 1.255 1.86 1.255 1.82 1.515 1.82 1.515 0.64 1.195 0.64 1.195 0.4 1.315 0.4 1.315 0.52 1.635 0.52 1.635 0.97 2.135 0.97 ;
      POLYGON 1.395 1.7 1.275 1.7 1.275 1 1.035 1 1.035 0.88 0.24 0.88 0.24 1.845 0.255 1.845 0.255 2.085 0.135 2.085 0.135 1.965 0.12 1.965 0.12 0.52 0.135 0.52 0.135 0.4 0.255 0.4 0.255 0.64 0.24 0.64 0.24 0.76 1.395 0.76 ;
  END
END MX2X1

MACRO SEDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX4 0 0 ;
  SIZE 13.63 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 0.63 1.515 1.99 ;
        RECT 0.555 1.025 1.515 1.145 ;
        RECT 0.555 0.885 0.8 1.145 ;
        RECT 0.555 0.63 0.675 1.99 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 1.03 8.395 1.44 ;
        RECT 8.135 1.15 8.395 1.38 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.77 1.14 9.005 1.46 ;
        RECT 8.77 1.135 8.92 1.46 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.18 11.005 1.41 ;
        RECT 10.845 1 10.965 1.41 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.485 1.21 12.865 1.4 ;
        RECT 12.485 1.21 12.745 1.425 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.005 0.97 13.125 1.21 ;
        RECT 12.775 0.94 13.035 1.09 ;
        RECT 11.845 0.97 13.125 1.09 ;
        RECT 11.725 1.28 11.965 1.4 ;
        RECT 11.845 0.97 11.965 1.4 ;
    END
  END E
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.63 0.18 ;
        RECT 12.845 -0.18 12.965 0.82 ;
        RECT 11.245 -0.18 11.365 0.64 ;
        RECT 8.525 0.51 8.765 0.63 ;
        RECT 8.525 -0.18 8.645 0.63 ;
        RECT 7.07 -0.18 7.19 0.73 ;
        RECT 4.655 0.49 4.895 0.61 ;
        RECT 4.775 -0.18 4.895 0.61 ;
        RECT 2.775 -0.18 2.895 0.68 ;
        RECT 1.815 -0.18 1.935 0.68 ;
        RECT 0.975 -0.18 1.095 0.68 ;
        RECT 0.135 -0.18 0.255 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.63 2.79 ;
        RECT 12.685 1.785 12.805 2.79 ;
        RECT 11.305 1.77 11.425 2.79 ;
        RECT 8.665 2.18 8.785 2.79 ;
        RECT 6.935 1.88 7.055 2.79 ;
        RECT 6.815 1.88 7.055 2 ;
        RECT 4.775 1.7 4.895 2.79 ;
        RECT 4.655 1.7 4.895 1.93 ;
        RECT 2.715 1.92 2.835 2.79 ;
        RECT 1.815 1.47 1.935 2.79 ;
        RECT 0.975 1.34 1.095 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.385 0.82 13.365 0.82 13.365 1.68 13.285 1.68 13.285 1.8 13.165 1.8 13.165 1.665 12.185 1.665 12.185 1.24 12.305 1.24 12.305 1.545 13.245 1.545 13.245 0.7 13.265 0.7 13.265 0.58 13.385 0.58 ;
      POLYGON 12.325 0.85 11.605 0.85 11.605 1.53 12.065 1.53 12.065 2.21 11.945 2.21 11.945 1.65 10.265 1.65 10.265 1.68 9.965 1.68 9.965 2.01 9.845 2.01 9.845 1.56 10.145 1.56 10.145 0.82 10.005 0.82 10.005 0.7 10.265 0.7 10.265 1.53 11.485 1.53 11.485 0.73 12.205 0.73 12.205 0.59 12.325 0.59 ;
      POLYGON 11.365 1.09 11.125 1.09 11.125 0.88 11.005 0.88 11.005 0.53 10.74 0.53 10.74 0.52 9.27 0.52 9.27 0.84 9.005 0.84 9.005 0.87 8.285 0.87 8.285 0.52 7.61 0.52 7.61 0.8 7.775 0.8 7.775 1.58 7.655 1.58 7.655 0.92 7.49 0.92 7.49 0.4 8.405 0.4 8.405 0.75 8.885 0.75 8.885 0.72 9.15 0.72 9.15 0.4 10.86 0.4 10.86 0.41 11.125 0.41 11.125 0.76 11.245 0.76 11.245 0.97 11.365 0.97 ;
      POLYGON 10.945 2.25 9.605 2.25 9.605 1.44 9.365 1.44 9.365 1.2 9.485 1.2 9.485 1.32 9.905 1.32 9.905 0.98 10.025 0.98 10.025 1.44 9.725 1.44 9.725 2.13 10.825 2.13 10.825 1.77 10.945 1.77 ;
      POLYGON 10.865 0.77 10.625 0.77 10.625 1.09 10.385 1.09 10.385 0.97 10.505 0.97 10.505 0.65 10.865 0.65 ;
      POLYGON 9.765 1.08 9.245 1.08 9.245 1.56 9.485 1.56 9.485 2.21 9.365 2.21 9.365 1.68 9.245 1.68 9.245 2.06 7.175 2.06 7.175 1.76 6.115 1.76 6.115 1.99 5.995 1.99 5.995 1.47 6.095 1.47 6.095 0.72 5.995 0.72 5.995 0.6 6.235 0.6 6.235 0.72 6.215 0.72 6.215 1.64 7.295 1.64 7.295 1.94 9.125 1.94 9.125 0.96 9.645 0.96 9.645 0.64 9.765 0.64 ;
      POLYGON 8.305 1.82 7.415 1.82 7.415 1.52 6.695 1.52 6.695 1.28 6.655 1.28 6.655 1 6.775 1 6.775 1.16 6.815 1.16 6.815 1.4 7.535 1.4 7.535 1.7 7.895 1.7 7.895 0.79 8.045 0.79 8.045 0.64 8.165 0.64 8.165 0.91 8.015 0.91 8.015 1.56 8.305 1.56 ;
      POLYGON 6.71 0.81 6.535 0.81 6.535 1.4 6.575 1.4 6.575 1.52 6.335 1.52 6.335 1.4 6.415 1.4 6.415 0.69 6.59 0.69 6.59 0.57 6.355 0.57 6.355 0.48 5.875 0.48 5.875 1.11 5.975 1.11 5.975 1.35 5.855 1.35 5.855 1.23 5.755 1.23 5.755 0.48 5.275 0.48 5.275 0.86 5.395 0.86 5.395 1.1 5.155 1.1 5.155 0.85 4.415 0.85 4.415 0.48 3.935 0.48 3.935 0.86 3.975 0.86 3.975 1.1 3.815 1.1 3.815 0.48 3.335 0.48 3.335 0.84 3.395 0.84 3.395 1.32 3.275 1.32 3.275 0.96 3.215 0.96 3.215 0.36 4.535 0.36 4.535 0.73 5.155 0.73 5.155 0.36 6.475 0.36 6.475 0.45 6.71 0.45 ;
      POLYGON 6.695 2.23 5.13 2.23 5.13 1.58 4.535 1.58 4.535 2.23 3.265 2.23 3.265 1.8 2.735 1.8 2.735 1.39 2.355 1.39 2.355 1.99 2.235 1.99 2.235 1.51 2.155 1.51 2.155 1.2 1.635 1.2 1.635 1.08 2.155 1.08 2.155 0.67 2.235 0.67 2.235 0.54 2.355 0.54 2.355 0.79 2.275 0.79 2.275 1.27 2.735 1.27 2.735 1.15 2.855 1.15 2.855 1.68 3.385 1.68 3.385 2.11 4.415 2.11 4.415 1.46 5.25 1.46 5.25 2.11 6.695 2.11 ;
      POLYGON 5.635 1.99 5.515 1.99 5.515 1.34 4.575 1.34 4.575 1.33 4.455 1.33 4.455 1.21 4.695 1.21 4.695 1.22 5.515 1.22 5.515 0.72 5.395 0.72 5.395 0.6 5.635 0.6 ;
      POLYGON 5.035 1.09 4.295 1.09 4.295 1.99 4.175 1.99 4.175 0.72 4.055 0.72 4.055 0.6 4.295 0.6 4.295 0.97 5.035 0.97 ;
      POLYGON 3.695 0.72 3.635 0.72 3.635 1.99 3.515 1.99 3.515 1.56 2.975 1.56 2.975 1.03 2.515 1.03 2.515 1.15 2.395 1.15 2.395 0.91 3.095 0.91 3.095 1.44 3.515 1.44 3.515 0.72 3.455 0.72 3.455 0.6 3.695 0.6 ;
  END
END SEDFFHQX4

MACRO OR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4XL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.02 1.675 1.455 ;
        RECT 1.535 1.02 1.66 1.48 ;
    END
  END A
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.51 1.63 ;
        RECT 0.36 1.175 0.48 1.66 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.125 0.82 1.54 ;
        RECT 0.7 1.105 0.82 1.54 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 1.33 1.16 1.66 ;
        RECT 0.94 1.175 1.09 1.51 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.055 2.44 1.175 ;
        RECT 2.32 0.66 2.44 1.175 ;
        RECT 2.1 1.055 2.25 1.435 ;
        RECT 2.1 1.055 2.22 1.96 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.9 -0.18 2.02 0.9 ;
        RECT 1.04 -0.18 1.16 0.38 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.68 1.84 1.8 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.98 1.72 1.4 1.72 1.4 1.9 0.16 1.9 0.16 1.78 1.28 1.78 1.28 0.9 0.56 0.9 0.56 0.66 0.68 0.66 0.68 0.78 1.48 0.78 1.48 0.66 1.6 0.66 1.6 0.9 1.4 0.9 1.4 1.6 1.86 1.6 1.86 1.38 1.98 1.38 ;
  END
END OR4XL

MACRO FILL8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL8 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
    END
  END VSS
END FILL8

MACRO EDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX8 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.03 0.51 1.485 ;
        RECT 0.36 1.03 0.48 1.515 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.255 11.085 1.465 ;
        RECT 10.745 1.23 11.005 1.465 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.035 0.99 11.405 1.11 ;
        RECT 10.505 0.97 11.295 1.09 ;
        RECT 11.035 0.94 11.295 1.11 ;
        RECT 10.725 0.41 10.845 1.09 ;
        RECT 10.025 0.41 10.845 0.53 ;
        RECT 10.025 0.41 10.145 1.01 ;
        RECT 10.005 0.89 10.125 1.46 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.045 0.8 8.045 0.92 ;
        RECT 7.925 0.68 8.045 0.92 ;
        RECT 7.625 1.45 7.865 1.59 ;
        RECT 5.045 1.45 7.865 1.57 ;
        RECT 6.965 0.68 7.085 0.92 ;
        RECT 6.785 1.45 7.025 1.59 ;
        RECT 5.885 1.45 6.125 1.59 ;
        RECT 6.005 0.68 6.125 0.92 ;
        RECT 5.58 1.175 5.73 1.57 ;
        RECT 5.61 0.8 5.73 1.57 ;
        RECT 5.045 1.45 5.285 1.59 ;
        RECT 5.045 0.68 5.165 0.92 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.065 -0.18 11.185 0.82 ;
        RECT 9.305 -0.18 9.425 0.64 ;
        RECT 8.405 0.46 8.645 0.58 ;
        RECT 8.525 -0.18 8.645 0.58 ;
        RECT 7.385 -0.18 7.625 0.32 ;
        RECT 6.425 -0.18 6.665 0.32 ;
        RECT 5.465 -0.18 5.705 0.32 ;
        RECT 4.565 -0.18 4.685 0.68 ;
        RECT 2.725 0.43 2.965 0.55 ;
        RECT 2.845 -0.18 2.965 0.55 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 11.005 1.825 11.125 2.79 ;
        RECT 9.305 2.1 9.545 2.22 ;
        RECT 9.305 2.1 9.425 2.79 ;
        RECT 8.345 2.1 8.585 2.22 ;
        RECT 8.345 2.1 8.465 2.79 ;
        RECT 7.205 1.95 7.445 2.07 ;
        RECT 7.205 1.95 7.325 2.79 ;
        RECT 6.305 1.95 6.545 2.075 ;
        RECT 6.305 1.95 6.425 2.79 ;
        RECT 5.465 1.95 5.705 2.075 ;
        RECT 5.465 1.95 5.585 2.79 ;
        RECT 4.625 1.95 4.865 2.075 ;
        RECT 4.625 1.95 4.745 2.79 ;
        RECT 2.725 1.75 2.845 2.79 ;
        RECT 0.555 1.635 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.645 1.705 11.605 1.705 11.605 1.825 11.485 1.825 11.485 1.705 10.505 1.705 10.505 1.24 10.625 1.24 10.625 1.585 11.525 1.585 11.525 0.82 11.485 0.82 11.485 0.58 11.605 0.58 11.605 0.7 11.645 0.7 ;
      POLYGON 10.605 0.77 10.485 0.77 10.485 0.85 10.385 0.85 10.385 2.21 10.265 2.21 10.265 1.98 8.265 1.98 8.265 1.83 4.41 1.83 4.41 2.17 4.145 2.17 4.145 2.23 2.965 2.23 2.965 1.63 2.555 1.63 2.555 2.23 1.545 2.23 1.545 1.59 1.425 1.59 1.425 0.72 1.305 0.72 1.305 0.6 1.545 0.6 1.545 1.47 1.665 1.47 1.665 2.11 2.435 2.11 2.435 1.51 3.085 1.51 3.085 2.11 4.025 2.11 4.025 2.05 4.29 2.05 4.29 1.71 8.385 1.71 8.385 1.86 10.265 1.86 10.265 0.73 10.365 0.73 10.365 0.65 10.605 0.65 ;
      POLYGON 10.025 1.74 9.765 1.74 9.765 1.62 9.065 1.62 9.065 1.74 8.825 1.74 8.825 1.62 8.885 1.62 8.885 1.33 7.065 1.33 7.065 1.13 7.305 1.13 7.305 1.21 8.885 1.21 8.885 0.59 9.005 0.59 9.005 0.76 9.665 0.76 9.665 0.65 9.905 0.65 9.905 0.77 9.785 0.77 9.785 0.88 9.005 0.88 9.005 1.5 9.885 1.5 9.885 1.62 10.025 1.62 ;
      POLYGON 8.765 1.09 8.525 1.09 8.525 0.82 8.165 0.82 8.165 0.56 4.925 0.56 4.925 0.92 4.485 0.92 4.485 1.59 4.17 1.59 4.17 1.65 4.165 1.65 4.165 1.93 3.925 1.93 3.925 1.53 4.05 1.53 4.05 1.47 4.365 1.47 4.365 0.92 3.925 0.92 3.925 0.54 4.045 0.54 4.045 0.8 4.805 0.8 4.805 0.44 8.285 0.44 8.285 0.7 8.645 0.7 8.645 0.97 8.765 0.97 ;
      POLYGON 4.245 1.35 4.125 1.35 4.125 1.16 3.685 1.16 3.685 1.12 3.565 1.12 3.565 0.88 3.685 0.88 3.685 0.48 3.205 0.48 3.205 0.79 2.385 0.79 2.385 1.12 2.245 1.12 2.245 0.88 2.265 0.88 2.265 0.48 1.785 0.48 1.785 0.84 1.805 0.84 1.805 1.35 1.685 1.35 1.685 0.96 1.665 0.96 1.665 0.48 1.135 0.48 1.135 1.635 1.095 1.635 1.095 1.755 0.975 1.755 0.975 1.515 1.015 1.515 1.015 0.67 0.975 0.67 0.975 0.36 2.605 0.36 2.605 0.67 3.085 0.67 3.085 0.36 3.805 0.36 3.805 1.04 4.245 1.04 ;
      POLYGON 3.565 0.72 3.445 0.72 3.445 1.99 3.325 1.99 3.325 1.39 2.745 1.39 2.745 1.15 2.865 1.15 2.865 1.27 3.325 1.27 3.325 0.6 3.565 0.6 ;
      POLYGON 3.205 1.15 3.085 1.15 3.085 1.03 2.625 1.03 2.625 1.36 2.125 1.36 2.125 1.99 2.005 1.99 2.005 0.72 1.905 0.72 1.905 0.6 2.145 0.6 2.145 0.72 2.125 0.72 2.125 1.24 2.505 1.24 2.505 0.91 3.205 0.91 ;
      POLYGON 0.895 0.95 0.655 0.95 0.655 0.91 0.24 0.91 0.24 1.635 0.255 1.635 0.255 1.875 0.135 1.875 0.135 1.755 0.12 1.755 0.12 0.67 0.135 0.67 0.135 0.43 0.255 0.43 0.255 0.79 0.895 0.79 ;
  END
END EDFFHQX8

MACRO AND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.415 1.295 ;
        RECT 0.295 1.055 0.415 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.465 1.09 1.82 ;
        RECT 0.815 1.465 1.09 1.61 ;
        RECT 0.815 1.25 0.935 1.61 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.485 1.435 1.605 1.83 ;
        RECT 1.35 1.435 1.605 1.555 ;
        RECT 1.23 1.175 1.47 1.435 ;
        RECT 1.35 0.53 1.47 1.555 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.93 -0.18 1.05 0.77 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.005 2.23 1.125 2.79 ;
        RECT 0.135 1.71 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.11 1.13 0.675 1.13 0.675 1.83 0.555 1.83 0.555 0.935 0.29 0.935 0.29 0.53 0.41 0.53 0.41 0.815 0.675 0.815 0.675 1.01 0.99 1.01 0.99 0.89 1.11 0.89 ;
  END
END AND2XL

MACRO CLKBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX3 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1 1.67 1.5 ;
        RECT 1.52 1 1.67 1.47 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.32 1.095 2.21 ;
        RECT 0.975 0.4 1.095 0.64 ;
        RECT 0.135 0.76 1.09 0.88 ;
        RECT 0.135 1.32 1.095 1.44 ;
        RECT 0.97 0.52 1.09 0.88 ;
        RECT 0.36 1.175 0.51 1.44 ;
        RECT 0.36 0.76 0.48 1.44 ;
        RECT 0.135 1.32 0.255 2.21 ;
        RECT 0.135 0.59 0.255 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.395 1.62 1.515 2.79 ;
        RECT 0.555 1.56 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 2.21 1.815 2.21 1.815 0.88 1.33 0.88 1.33 1.17 1.21 1.17 1.21 0.76 1.815 0.76 1.815 0.59 1.935 0.59 ;
  END
END CLKBUFX3

MACRO DFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRXL 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.965 1.27 2.085 1.51 ;
        RECT 1.84 1.39 2.085 1.51 ;
        RECT 1.81 1.465 1.96 1.725 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.74 1.025 7.095 1.16 ;
        RECT 6.74 0.885 6.89 1.18 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.335 0.735 7.455 1.24 ;
        RECT 7.03 0.735 7.455 0.855 ;
        RECT 7.03 0.595 7.18 0.855 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 1.31 1.485 1.83 ;
        RECT 1.365 0.67 1.485 0.91 ;
        RECT 1.23 1.175 1.445 1.435 ;
        RECT 1.325 0.79 1.445 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 6.865 -0.18 6.985 0.38 ;
        RECT 4.73 -0.18 4.97 0.32 ;
        RECT 3.135 -0.18 3.255 0.9 ;
        RECT 1.785 -0.18 1.905 0.39 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.575 1.98 7.695 2.79 ;
        RECT 6.835 1.98 6.955 2.79 ;
        RECT 4.715 2.16 4.955 2.28 ;
        RECT 4.715 2.16 4.835 2.79 ;
        RECT 3.015 2.16 3.255 2.28 ;
        RECT 3.015 2.16 3.135 2.79 ;
        RECT 1.725 2.23 1.845 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.695 1.48 7.315 1.48 7.315 1.76 6.015 1.76 6.015 1.86 5.895 1.86 5.895 1.62 6.055 1.62 6.055 0.9 5.995 0.9 5.995 0.66 6.115 0.66 6.115 0.78 6.175 0.78 6.175 1.64 7.195 1.64 7.195 1.36 7.575 1.36 7.575 0.66 7.695 0.66 ;
      POLYGON 6.535 1.52 6.295 1.52 6.295 1.4 6.385 1.4 6.385 0.66 6.285 0.66 6.285 0.54 5.875 0.54 5.875 1.36 5.935 1.36 5.935 1.48 5.695 1.48 5.695 1.36 5.755 1.36 5.755 0.54 5.21 0.54 5.21 0.56 4.175 0.56 4.175 1 4.315 1 4.315 1.24 4.055 1.24 4.055 1.14 3.755 1.14 3.755 1.54 3.635 1.54 3.635 1.02 4.055 1.02 4.055 0.44 5.09 0.44 5.09 0.42 5.235 0.42 5.235 0.38 5.475 0.38 5.475 0.42 6.405 0.42 6.405 0.54 6.505 0.54 6.505 1.4 6.535 1.4 ;
      POLYGON 5.635 0.84 5.575 0.84 5.575 1.62 5.595 1.62 5.595 1.86 5.475 1.86 5.475 1.74 5.455 1.74 5.455 1.48 4.675 1.48 4.675 1.36 5.455 1.36 5.455 0.84 5.395 0.84 5.395 0.72 5.635 0.72 ;
      POLYGON 5.515 2.24 5.275 2.24 5.275 2.1 5.175 2.1 5.175 2.04 4.235 2.04 4.235 2.24 3.995 2.24 3.995 2.04 2.205 2.04 2.205 1.68 2.265 1.68 2.265 0.67 2.385 0.67 2.385 1.8 2.325 1.8 2.325 1.92 5.295 1.92 5.295 1.98 5.395 1.98 5.395 2.12 5.515 2.12 ;
      POLYGON 5.135 1.16 4.555 1.16 4.555 1.8 4.235 1.8 4.235 1.68 4.435 1.68 4.435 0.84 4.295 0.84 4.295 0.72 4.555 0.72 4.555 1.04 5.135 1.04 ;
      POLYGON 3.955 1.8 3.715 1.8 3.715 1.78 3.395 1.78 3.395 1.5 2.915 1.5 2.915 1.46 2.755 1.46 2.755 1.34 3.035 1.34 3.035 1.38 3.395 1.38 3.395 0.78 3.815 0.78 3.815 0.66 3.935 0.66 3.935 0.9 3.515 0.9 3.515 1.66 3.835 1.66 3.835 1.68 3.955 1.68 ;
      POLYGON 3.275 1.26 3.155 1.26 3.155 1.22 2.635 1.22 2.635 1.68 2.775 1.68 2.775 1.8 2.515 1.8 2.515 0.78 2.655 0.78 2.655 0.66 2.555 0.66 2.555 0.55 2.145 0.55 2.145 1.15 1.805 1.15 1.805 1.19 1.565 1.19 1.565 1.03 2.025 1.03 2.025 0.43 2.675 0.43 2.675 0.54 2.775 0.54 2.775 0.9 2.635 0.9 2.635 1.1 3.155 1.1 3.155 1.02 3.275 1.02 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFTRXL

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.98 0.355 1.22 ;
        RECT 0.07 0.98 0.355 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.215 1.145 1.38 ;
        RECT 0.775 1.2 0.895 1.475 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.505 0.885 1.67 1.145 ;
        RECT 1.355 1.36 1.625 1.48 ;
        RECT 1.505 0.72 1.625 1.48 ;
        RECT 1.355 0.72 1.625 0.84 ;
        RECT 1.355 1.36 1.475 2.21 ;
        RECT 1.355 0.6 1.475 0.84 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 1.775 -0.18 1.895 0.73 ;
        RECT 0.875 0.72 1.115 0.84 ;
        RECT 0.875 -0.18 0.995 0.84 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 1.56 1.895 2.79 ;
        RECT 0.935 1.595 1.055 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.385 1.24 1.265 1.24 1.265 1.08 0.635 1.08 0.635 1.46 0.415 1.46 0.415 1.74 0.175 1.74 0.175 1.62 0.295 1.62 0.295 1.34 0.515 1.34 0.515 0.66 0.635 0.66 0.635 0.96 1.385 0.96 ;
  END
END OR2X2

MACRO DLY2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X4 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.6 1.515 2.21 ;
        RECT 1.215 0.52 1.515 0.64 ;
        RECT 1.395 0.4 1.515 0.64 ;
        RECT 1.215 1.6 1.515 1.72 ;
        RECT 1.215 0.52 1.335 1.72 ;
        RECT 0.555 0.885 1.335 1.005 ;
        RECT 0.555 0.885 0.8 1.145 ;
        RECT 0.555 0.59 0.675 2.21 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 0.77 3.7 1.145 ;
        RECT 3.505 1.02 3.625 1.4 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.24 1.48 6.66 1.72 ;
        RECT 6.54 0.98 6.66 1.72 ;
        RECT 6.365 0.98 6.66 1.1 ;
        RECT 6.365 -0.18 6.485 1.1 ;
        RECT 5.765 0.68 6.005 0.8 ;
        RECT 5.765 -0.18 5.885 0.8 ;
        RECT 4.205 1.3 4.485 1.42 ;
        RECT 4.365 -0.18 4.485 1.42 ;
        RECT 3.645 -0.18 3.885 0.32 ;
        RECT 2.455 1.1 2.735 1.22 ;
        RECT 2.615 -0.18 2.735 1.22 ;
        RECT 1.815 -0.18 1.935 0.64 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 5.22 1.22 6.42 1.34 ;
        RECT 5.22 1.84 5.58 2.15 ;
        RECT 5.22 1.84 5.46 2.79 ;
        RECT 5.22 1.06 5.34 2.79 ;
        RECT 5.085 1.06 5.34 1.18 ;
        RECT 3.725 2.18 3.845 2.79 ;
        RECT 2.255 0.76 2.495 0.9 ;
        RECT 1.455 0.76 2.495 0.88 ;
        RECT 1.635 1.82 1.995 2.15 ;
        RECT 1.635 1.82 1.875 2.79 ;
        RECT 1.635 1.36 1.755 2.79 ;
        RECT 1.455 1.36 1.755 1.48 ;
        RECT 1.455 0.76 1.575 1.48 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.9 1.98 6.32 1.98 6.32 1.96 6 1.96 6 1.72 5.66 1.72 5.66 1.46 5.78 1.46 5.78 1.6 6.12 1.6 6.12 1.84 6.78 1.84 6.78 0.86 6.605 0.86 6.605 0.62 6.725 0.62 6.725 0.74 6.9 0.74 ;
      POLYGON 6.245 1.04 5.525 1.04 5.525 0.62 4.99 0.62 4.99 0.68 4.725 0.68 4.725 1.7 4.545 1.7 4.545 1.82 4.425 1.82 4.425 1.58 4.605 1.58 4.605 0.56 4.87 0.56 4.87 0.5 5.645 0.5 5.645 0.92 6.125 0.92 6.125 0.48 6.005 0.48 6.005 0.36 6.245 0.36 ;
      POLYGON 5.405 0.86 5.285 0.86 5.285 0.94 4.965 0.94 4.965 1.56 5.1 1.56 5.1 2.21 4.98 2.21 4.98 2.06 3.56 2.06 3.56 2.22 2.115 2.22 2.115 1.7 1.875 1.7 1.875 1.24 1.695 1.24 1.695 1 1.815 1 1.815 1.12 1.995 1.12 1.995 1.58 2.235 1.58 2.235 2.1 3.44 2.1 3.44 1.94 4.845 1.94 4.845 0.82 5.165 0.82 5.165 0.74 5.405 0.74 ;
      POLYGON 4.245 0.54 4.125 0.54 4.125 0.56 2.975 0.56 2.975 1.46 2.835 1.46 2.835 1.74 2.595 1.74 2.595 1.62 2.715 1.62 2.715 1.34 2.855 1.34 2.855 0.4 2.975 0.4 2.975 0.44 4.005 0.44 4.005 0.42 4.245 0.42 ;
      POLYGON 3.365 1.82 3.32 1.82 3.32 1.98 2.355 1.98 2.355 1.46 2.115 1.46 2.115 1.22 2.235 1.22 2.235 1.34 2.475 1.34 2.475 1.86 3.2 1.86 3.2 1.7 3.245 1.7 3.245 0.68 3.365 0.68 ;
  END
END DLY2X4

MACRO MXI4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X2 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.42 1.145 4.57 1.435 ;
        RECT 4.31 1.14 4.43 1.42 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 1.23 7.815 1.38 ;
        RECT 7.555 1.14 7.795 1.38 ;
        RECT 7.475 1.38 7.63 1.5 ;
        RECT 7.21 1.555 7.595 1.675 ;
        RECT 7.475 1.38 7.595 1.675 ;
        RECT 7.51 1.26 7.595 1.675 ;
        RECT 4.93 1.96 7.33 2.08 ;
        RECT 7.21 1.555 7.33 2.08 ;
        RECT 5.01 1.24 5.13 1.48 ;
        RECT 4.93 1.36 5.05 2.08 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.5 1.03 1.63 ;
        RECT 0.65 1.465 0.8 1.75 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.54 2.425 1.78 ;
        RECT 2.045 1.52 2.305 1.78 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3288 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.8267 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 1.16 1.33 1.4 ;
        RECT 0.36 1.225 1.33 1.345 ;
        RECT 0.41 1.225 0.53 1.465 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.54 2.93 1.77 ;
        RECT 2.625 1.52 2.885 1.77 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.97 1.175 7.18 1.435 ;
        RECT 6.97 0.74 7.09 1.84 ;
        RECT 6.85 0.74 7.09 0.86 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.45 -0.18 7.57 0.78 ;
        RECT 6.13 0.6 6.37 0.72 ;
        RECT 6.13 -0.18 6.25 0.72 ;
        RECT 4.33 -0.18 4.45 0.78 ;
        RECT 2.49 -0.18 2.61 0.68 ;
        RECT 0.65 -0.18 0.77 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.45 2.06 7.57 2.79 ;
        RECT 6.49 2.2 6.61 2.79 ;
        RECT 4.39 2.28 4.63 2.79 ;
        RECT 2.49 2.14 2.61 2.79 ;
        RECT 0.59 1.96 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.055 1.62 7.75 1.62 7.75 1.5 7.935 1.5 7.935 1.02 7.21 1.02 7.21 0.62 6.61 0.62 6.61 1.6 5.41 1.6 5.41 1.12 4.93 1.12 4.93 1.06 4.81 1.06 4.81 0.94 5.05 0.94 5.05 1 5.53 1 5.53 1.48 6.49 1.48 6.49 0.5 7.33 0.5 7.33 0.9 7.93 0.9 7.93 0.66 8.05 0.66 8.05 0.78 8.055 0.78 ;
      POLYGON 6.85 1.84 5.17 1.84 5.17 1.6 5.29 1.6 5.29 1.72 6.73 1.72 6.73 1.18 6.85 1.18 ;
      POLYGON 6.37 1.36 5.65 1.36 5.65 0.88 5.17 0.88 5.17 0.72 4.97 0.72 4.97 0.6 5.29 0.6 5.29 0.76 5.77 0.76 5.77 1.24 6.37 1.24 ;
      POLYGON 6.13 1.04 5.89 1.04 5.89 0.48 4.69 0.48 4.69 1.02 4.19 1.02 4.19 1.92 3.81 1.92 3.81 2 3.57 2 3.57 1.88 3.69 1.88 3.69 1.8 4.07 1.8 4.07 0.88 3.63 0.88 3.63 0.62 3.75 0.62 3.75 0.76 4.19 0.76 4.19 0.9 4.57 0.9 4.57 0.36 6.01 0.36 6.01 0.92 6.13 0.92 ;
      POLYGON 4.81 2.16 4.05 2.16 4.05 2.24 3.305 2.24 3.305 2.02 1.57 2.02 1.57 2.08 1.45 2.08 1.45 0.62 1.57 0.62 1.57 1.9 3.425 1.9 3.425 2.12 3.93 2.12 3.93 2.04 4.69 2.04 4.69 1.24 4.81 1.24 ;
      POLYGON 3.95 1.12 3.83 1.12 3.83 1.4 3.19 1.4 3.19 1.72 3.07 1.72 3.07 1.4 1.93 1.4 1.93 1.16 2.05 1.16 2.05 1.28 3.71 1.28 3.71 1 3.95 1 ;
      POLYGON 3.95 1.68 3.71 1.68 3.71 1.64 3.35 1.64 3.35 1.52 3.83 1.52 3.83 1.56 3.95 1.56 ;
      RECT 2.99 1.04 3.59 1.16 ;
      POLYGON 3.23 0.48 3.11 0.48 3.11 0.92 2.195 0.92 2.195 0.5 1.81 0.5 1.81 1.76 1.69 1.76 1.69 0.5 1.015 0.5 1.015 1.04 0.24 1.04 0.24 1.555 0.29 1.555 0.29 2.08 0.17 2.08 0.17 1.675 0.12 1.675 0.12 0.8 0.17 0.8 0.17 0.68 0.29 0.68 0.29 0.92 0.895 0.92 0.895 0.38 1.16 0.38 1.16 0.36 1.4 0.36 1.4 0.38 2.315 0.38 2.315 0.8 2.99 0.8 2.99 0.36 3.23 0.36 ;
  END
END MXI4X2

MACRO TLATNXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNXL 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.72 1.04 0.84 1.42 ;
        RECT 0.65 1.065 0.8 1.435 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.275 3.41 1.725 ;
        RECT 3.29 1.25 3.41 1.725 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.93 1.585 4.05 2.09 ;
        RECT 3.84 1.345 3.99 1.725 ;
        RECT 3.81 0.64 3.93 1.465 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.16 1.435 5.28 1.675 ;
        RECT 5 1.175 5.16 1.435 ;
        RECT 5.04 0.575 5.16 1.555 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.62 -0.18 4.74 0.815 ;
        RECT 3.33 -0.18 3.45 0.88 ;
        RECT 2.04 -0.18 2.16 0.64 ;
        RECT 0.65 -0.18 0.77 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.74 1.555 4.86 2.79 ;
        RECT 3.51 1.97 3.63 2.79 ;
        RECT 2.3 2.08 2.42 2.79 ;
        RECT 0.615 2.08 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.88 1.075 4.44 1.075 4.44 1.675 4.32 1.675 4.32 0.955 4.2 0.955 4.2 0.575 4.32 0.575 4.32 0.835 4.44 0.835 4.44 0.955 4.88 0.955 ;
      POLYGON 3.81 0.48 3.69 0.48 3.69 1.12 3.09 1.12 3.09 0.52 2.73 0.52 2.73 1.48 2.9 1.48 2.9 1.72 2.78 1.72 2.78 1.6 2.61 1.6 2.61 1.24 2.27 1.24 2.27 1.36 2.15 1.36 2.15 1.12 2.61 1.12 2.61 0.64 2.46 0.64 2.46 0.4 3.21 0.4 3.21 1 3.57 1 3.57 0.36 3.81 0.36 ;
      POLYGON 3.21 2.11 3.09 2.11 3.09 1.99 3.02 1.99 3.02 1.965 2.56 1.965 2.56 1.96 1.36 1.96 1.36 0.92 0.53 0.92 0.53 0.98 0.41 0.98 0.41 0.74 0.53 0.74 0.53 0.8 1.48 0.8 1.48 1.22 1.67 1.22 1.67 1.1 1.79 1.1 1.79 1.34 1.48 1.34 1.48 1.84 2.68 1.84 2.68 1.845 3.02 1.845 3.02 1.36 2.85 1.36 2.85 0.64 2.97 0.64 2.97 1.24 3.14 1.24 3.14 1.845 3.21 1.845 ;
      POLYGON 2.49 1 2.37 1 2.37 0.98 2.03 0.98 2.03 1.58 1.72 1.58 1.72 1.7 1.6 1.7 1.6 1.46 1.91 1.46 1.91 0.98 1.6 0.98 1.6 0.68 1.29 0.68 1.29 0.4 1.41 0.4 1.41 0.56 1.72 0.56 1.72 0.86 2.37 0.86 2.37 0.76 2.49 0.76 ;
      POLYGON 1.24 1.3 1.12 1.3 1.12 1.675 0.255 1.675 0.255 1.795 0.135 1.795 0.135 1.555 0.17 1.555 0.17 0.4 0.29 0.4 0.29 1.555 1 1.555 1 1.18 1.24 1.18 ;
  END
END TLATNXL

MACRO DFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX2 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 1.345 0.53 1.8 ;
        RECT 0.36 1.29 0.51 1.725 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 1.165 4.625 1.38 ;
        RECT 4.465 1 4.585 1.38 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.03 5.15 1.435 ;
        RECT 4.985 1 5.105 1.41 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.46 0.87 1.78 ;
        RECT 0.65 1.455 0.8 1.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.565 1.465 9.79 1.725 ;
        RECT 9.565 1.34 9.76 1.725 ;
        RECT 9.62 0.59 9.74 1.725 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 1.465 10.66 1.725 ;
        RECT 10.48 1.45 10.645 1.57 ;
        RECT 10.48 0.71 10.6 1.57 ;
        RECT 10.46 0.59 10.58 0.83 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.88 -0.18 11 0.64 ;
        RECT 10.04 -0.18 10.16 0.64 ;
        RECT 9.2 -0.18 9.32 0.73 ;
        RECT 7.07 -0.18 7.19 0.78 ;
        RECT 4.605 0.48 4.845 0.64 ;
        RECT 4.605 -0.18 4.725 0.64 ;
        RECT 2.15 -0.18 2.39 0.32 ;
        RECT 0.67 -0.18 0.79 0.86 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 11.005 2.085 11.125 2.79 ;
        RECT 10.045 2.085 10.165 2.79 ;
        RECT 9.085 1.86 9.205 2.79 ;
        RECT 7.97 1.87 8.31 1.99 ;
        RECT 8.19 1.63 8.31 1.99 ;
        RECT 7.97 1.87 8.09 2.79 ;
        RECT 7.13 1.86 7.25 2.79 ;
        RECT 4.19 2.275 4.43 2.79 ;
        RECT 3.005 2.1 3.125 2.79 ;
        RECT 2.19 2.1 2.31 2.79 ;
        RECT 0.59 1.92 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.465 1.58 11.345 1.58 11.345 0.88 10.84 0.88 10.84 1.17 10.72 1.17 10.72 0.76 11.3 0.76 11.3 0.4 11.42 0.4 11.42 0.76 11.465 0.76 ;
      POLYGON 11.16 1.965 9.325 1.965 9.325 1.74 8.725 1.74 8.725 2.25 8.21 2.25 8.21 2.13 8.605 2.13 8.605 1.62 9.305 1.62 9.305 1.01 8.78 1.01 8.78 0.59 8.9 0.59 8.9 0.89 9.425 0.89 9.425 1.62 9.445 1.62 9.445 1.845 9.91 1.845 9.91 1.26 9.9 1.26 9.9 1.02 10.03 1.02 10.03 1.845 11.04 1.845 11.04 1 11.16 1 ;
      POLYGON 8.885 1.5 6.32 1.5 6.32 1.77 6.2 1.77 6.2 0.67 6.32 0.67 6.32 1.38 8.765 1.38 8.765 1.13 8.885 1.13 ;
      POLYGON 8.51 1.02 7.6 1.02 7.6 0.84 7.55 0.84 7.55 0.6 7.67 0.6 7.67 0.72 7.72 0.72 7.72 0.9 8.39 0.9 8.39 0.6 8.51 0.6 ;
      POLYGON 8.23 1.26 6.44 1.26 6.44 0.55 5.265 0.55 5.265 0.76 5.39 0.76 5.39 1.41 5.51 1.41 5.51 1.53 5.27 1.53 5.27 0.88 4.305 0.88 4.305 0.48 4.065 0.48 4.065 0.36 4.425 0.36 4.425 0.76 4.965 0.76 4.965 0.64 5.145 0.64 5.145 0.43 6.56 0.43 6.56 1.14 8.23 1.14 ;
      POLYGON 8.15 0.78 7.91 0.78 7.91 0.66 7.84 0.66 7.84 0.48 7.43 0.48 7.43 1.02 6.68 1.02 6.68 0.67 6.8 0.67 6.8 0.9 7.31 0.9 7.31 0.36 7.96 0.36 7.96 0.54 8.03 0.54 8.03 0.66 8.15 0.66 ;
      POLYGON 7.67 1.98 7.55 1.98 7.55 1.86 7.37 1.86 7.37 1.74 6.56 1.74 6.56 1.62 7.49 1.62 7.49 1.74 7.67 1.74 ;
      POLYGON 6.52 2.15 6.22 2.15 6.22 2.01 4.79 2.01 4.79 1.915 3.885 1.915 3.885 1.36 2.81 1.36 2.81 1.24 4.005 1.24 4.005 1.795 4.91 1.795 4.91 1.89 5.96 1.89 5.96 1.23 5.9 1.23 5.9 0.99 6.02 0.99 6.02 1.11 6.08 1.11 6.08 1.89 6.34 1.89 6.34 2.03 6.52 2.03 ;
      POLYGON 6.1 2.25 4.55 2.25 4.55 2.155 3.645 2.155 3.645 2.01 3.485 2.01 3.485 1.74 2.55 1.74 2.55 1.44 1.57 1.44 1.57 1.32 2.57 1.32 2.57 0.92 2.55 0.92 2.55 0.68 2.67 0.68 2.67 0.8 2.69 0.8 2.69 1.62 3.605 1.62 3.605 1.89 3.765 1.89 3.765 2.035 4.67 2.035 4.67 2.13 6.1 2.13 ;
      POLYGON 5.84 1.77 5.03 1.77 5.03 1.675 4.125 1.675 4.125 1.12 2.925 1.12 2.925 0.56 1.91 0.56 1.91 0.48 1.79 0.48 1.79 0.36 2.03 0.36 2.03 0.44 3.045 0.44 3.045 1 3.585 1 3.585 0.64 3.705 0.64 3.705 1 4.245 1 4.245 1.5 4.365 1.5 4.365 1.555 5.15 1.555 5.15 1.65 5.66 1.65 5.66 0.67 5.78 0.67 5.78 1.53 5.84 1.53 ;
      POLYGON 4.185 0.82 3.825 0.82 3.825 0.52 3.465 0.52 3.465 0.64 3.285 0.64 3.285 0.88 3.165 0.88 3.165 0.52 3.345 0.52 3.345 0.4 3.945 0.4 3.945 0.7 4.185 0.7 ;
      POLYGON 3.525 2.25 3.245 2.25 3.245 1.98 1.45 1.98 1.45 2.04 1.33 2.04 1.33 1.36 1.31 1.36 1.31 0.62 1.43 0.62 1.43 1.24 1.45 1.24 1.45 1.86 3.365 1.86 3.365 2.13 3.525 2.13 ;
      POLYGON 2.45 1.18 1.57 1.18 1.57 0.94 1.55 0.94 1.55 0.5 1.19 0.5 1.19 1.48 1.21 1.48 1.21 1.72 1.07 1.72 1.07 1.17 0.24 1.17 0.24 1.845 0.29 1.845 0.29 2.085 0.17 2.085 0.17 1.965 0.12 1.965 0.12 0.74 0.25 0.74 0.25 0.62 0.37 0.62 0.37 0.86 0.24 0.86 0.24 1.05 1.07 1.05 1.07 0.38 1.67 0.38 1.67 0.82 1.69 0.82 1.69 1 1.81 1 1.81 1.06 2.45 1.06 ;
  END
END DFFNSRX2

MACRO OR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X4 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 0.51 1.45 ;
        RECT 0.36 1 0.48 1.475 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1 0.87 1.345 ;
        RECT 0.65 1.09 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.37 1.38 1.725 ;
        RECT 1.23 1.23 1.35 1.725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.885 3.12 1.145 ;
        RECT 2.71 0.885 3.12 1.005 ;
        RECT 2.57 1.56 2.83 1.68 ;
        RECT 2.71 0.71 2.83 1.68 ;
        RECT 2.67 0.59 2.79 0.83 ;
        RECT 1.73 1.32 2.83 1.44 ;
        RECT 2.57 1.56 2.69 2.21 ;
        RECT 1.89 0.71 2.83 0.83 ;
        RECT 1.77 0.65 2.01 0.77 ;
        RECT 1.73 1.32 1.85 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 3.09 -0.18 3.21 0.64 ;
        RECT 2.19 0.46 2.43 0.58 ;
        RECT 2.19 -0.18 2.31 0.58 ;
        RECT 1.41 -0.18 1.53 0.64 ;
        RECT 0.57 -0.18 0.69 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.99 1.56 3.11 2.79 ;
        RECT 2.15 1.56 2.27 2.79 ;
        RECT 1.31 1.845 1.43 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.59 1.11 1.11 1.11 1.11 1.715 0.39 1.715 0.39 2.21 0.27 2.21 0.27 1.595 0.99 1.595 0.99 0.88 0.15 0.88 0.15 0.59 0.27 0.59 0.27 0.76 0.99 0.76 0.99 0.59 1.11 0.59 1.11 0.99 2.59 0.99 ;
  END
END OR3X4

MACRO XOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2XL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.835 1.29 0.955 1.53 ;
        RECT 0.68 1.41 0.955 1.53 ;
        RECT 0.65 1.465 0.8 1.725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.415 1.27 2.655 1.39 ;
        RECT 1.335 1.17 2.535 1.29 ;
        RECT 1.855 1.09 2.095 1.29 ;
        RECT 1.755 1.17 2.015 1.38 ;
        RECT 1.335 1.17 1.455 1.55 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.55 0.255 1.87 ;
        RECT 0.07 1.465 0.255 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.355 0.61 2.595 0.73 ;
        RECT 2.355 -0.18 2.475 0.73 ;
        RECT 0.495 0.61 0.735 0.73 ;
        RECT 0.495 -0.18 0.615 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.215 1.75 2.335 2.79 ;
        RECT 0.615 2.23 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.955 0.79 2.895 0.79 2.895 1.75 2.755 1.75 2.755 1.87 2.635 1.87 2.635 1.63 1.895 1.63 1.895 2.25 1.655 2.25 1.655 2.13 1.775 2.13 1.775 1.51 2.775 1.51 2.775 0.67 2.835 0.67 2.835 0.55 2.955 0.55 ;
      POLYGON 2.455 1.05 2.215 1.05 2.215 0.97 1.215 0.97 1.215 1.87 1.095 1.87 1.095 0.61 1.335 0.61 1.335 0.73 1.215 0.73 1.215 0.85 2.335 0.85 2.335 0.93 2.455 0.93 ;
      POLYGON 1.955 0.73 1.715 0.73 1.715 0.49 0.975 0.49 0.975 1.17 0.53 1.17 0.53 1.845 0.74 1.845 0.74 1.99 1.415 1.99 1.415 1.87 1.515 1.87 1.515 1.75 1.635 1.75 1.635 1.99 1.535 1.99 1.535 2.11 0.62 2.11 0.62 1.965 0.41 1.965 0.41 0.95 0.53 0.95 0.53 1.05 0.855 1.05 0.855 0.37 1.835 0.37 1.835 0.61 1.955 0.61 ;
  END
END XOR2XL

MACRO DFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRXL 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 0.92 7.525 1.19 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.22 2.015 1.45 ;
        RECT 1.815 1.18 1.935 1.59 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3384 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.82 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.15 3.215 1.38 ;
        RECT 2.915 1.15 3.175 1.405 ;
    END
  END RN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1584 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 0.7 1.485 0.82 ;
        RECT 1.365 0.58 1.485 0.82 ;
        RECT 1.215 1.465 1.38 1.725 ;
        RECT 1.215 0.7 1.335 2.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.265 0.68 7.505 0.8 ;
        RECT 7.385 -0.18 7.505 0.8 ;
        RECT 5.375 0.47 5.615 0.59 ;
        RECT 5.495 -0.18 5.615 0.59 ;
        RECT 3.315 -0.18 3.435 0.75 ;
        RECT 1.785 -0.18 1.905 0.82 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.665 2.11 7.785 2.79 ;
        RECT 6.065 2.15 6.185 2.79 ;
        RECT 5.255 2.29 5.495 2.79 ;
        RECT 3.315 2.29 3.555 2.79 ;
        RECT 2.445 2.15 2.565 2.79 ;
        RECT 1.695 2.23 1.815 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.325 1.75 8.085 1.75 8.085 1.43 7.225 1.43 7.225 1.55 7.105 1.55 7.105 1.43 7.025 1.43 7.025 0.5 5.855 0.5 5.855 0.83 5.135 0.83 5.135 0.48 4.655 0.48 4.655 1.06 3.995 1.06 3.995 1.41 3.875 1.41 3.875 0.94 4.535 0.94 4.535 0.36 5.255 0.36 5.255 0.71 5.735 0.71 5.735 0.38 6.235 0.38 6.235 0.36 6.475 0.36 6.475 0.38 7.145 0.38 7.145 1.31 7.825 1.31 7.825 0.62 7.945 0.62 7.945 1.31 8.205 1.31 8.205 1.63 8.325 1.63 ;
      POLYGON 8.125 2.25 8.005 2.25 8.005 1.99 7.33 1.99 7.33 2.15 6.92 2.15 6.92 2.25 6.68 2.25 6.68 2.15 6.305 2.15 6.305 2.03 5.935 2.03 5.935 1.93 2.175 1.93 2.175 1.95 2.055 1.95 2.055 1.71 2.265 1.71 2.265 0.6 2.385 0.6 2.385 1.81 4.535 1.81 4.535 1.33 4.755 1.33 4.755 1.19 4.875 1.19 4.875 1.45 4.655 1.45 4.655 1.81 6.055 1.81 6.055 1.91 6.425 1.91 6.425 2.03 7.21 2.03 7.21 1.87 8.125 1.87 ;
      POLYGON 7.085 1.91 6.965 1.91 6.965 1.79 6.785 1.79 6.785 1.37 5.235 1.37 5.235 1.25 6.545 1.25 6.545 0.62 6.665 0.62 6.665 1.25 6.905 1.25 6.905 1.67 7.085 1.67 ;
      POLYGON 6.665 1.87 6.545 1.87 6.545 1.69 5.735 1.69 5.735 1.57 6.665 1.57 ;
      POLYGON 6.225 1.13 5.115 1.13 5.115 1.69 4.775 1.69 4.775 1.57 4.995 1.57 4.995 1.07 4.775 1.07 4.775 0.6 5.015 0.6 5.015 0.95 5.115 0.95 5.115 1.01 6.225 1.01 ;
      RECT 2.995 2.05 5.815 2.17 ;
      POLYGON 4.415 0.72 3.755 0.72 3.755 1.53 4.095 1.53 4.095 1.57 4.215 1.57 4.215 1.69 3.975 1.69 3.975 1.65 3.635 1.65 3.635 1.03 2.745 1.03 2.745 0.91 3.635 0.91 3.635 0.6 4.415 0.6 ;
      POLYGON 3.515 1.645 3.075 1.645 3.075 1.69 2.835 1.69 2.835 1.645 2.505 1.645 2.505 0.63 2.675 0.63 2.675 0.48 2.145 0.48 2.145 1.06 1.695 1.06 1.695 1.1 1.455 1.1 1.455 0.94 2.025 0.94 2.025 0.36 2.795 0.36 2.795 0.75 2.625 0.75 2.625 1.525 3.395 1.525 3.395 1.19 3.515 1.19 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFRXL

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 1.45 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 0.595 0.8 1.2 ;
        RECT 0.65 0.595 0.8 1.02 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.825 0.51 1.2 ;
        RECT 0.36 0.825 0.48 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3284 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 1.175 1.09 1.435 ;
        RECT 0.62 1.32 1.04 1.44 ;
        RECT 0.92 0.62 1.04 1.44 ;
        RECT 0.62 1.32 0.74 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.45 0.18 ;
        RECT 0.2 -0.18 0.32 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.45 2.79 ;
        RECT 1.04 1.56 1.16 2.79 ;
        RECT 0.2 1.56 0.32 2.79 ;
    END
  END VDD
END NAND2X1

MACRO FILL16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL16 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
    END
  END VSS
END FILL16

MACRO CLKBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX6 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 1.39 2.01 2.21 ;
        RECT 0.15 0.91 2.01 1.03 ;
        RECT 1.89 0.4 2.01 1.03 ;
        RECT 0.21 1.39 2.01 1.51 ;
        RECT 1.05 1.39 1.17 2.21 ;
        RECT 0.99 0.4 1.11 1.03 ;
        RECT 0.36 1.175 0.51 1.51 ;
        RECT 0.36 0.91 0.48 1.51 ;
        RECT 0.21 1.39 0.33 2.21 ;
        RECT 0.15 0.4 0.27 1.03 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.825 3.12 1.285 ;
        RECT 2.97 0.825 3.09 1.31 ;
    END
  END A
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 3.15 1.43 3.27 2.79 ;
        RECT 2.31 1.43 2.43 2.79 ;
        RECT 1.47 1.63 1.59 2.79 ;
        RECT 0.63 1.63 0.75 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 3.15 -0.18 3.27 0.705 ;
        RECT 2.31 -0.18 2.43 0.895 ;
        RECT 1.41 -0.18 1.53 0.79 ;
        RECT 0.57 -0.18 0.69 0.79 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.85 2.08 2.73 2.08 2.73 1.27 0.77 1.27 0.77 1.15 2.73 1.15 2.73 0.655 2.85 0.655 ;
  END
END CLKBUFX6

MACRO AOI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222XL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 0.915 1.145 1.105 ;
        RECT 0.705 0.88 1.005 1.035 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.37 0.71 2.54 1.145 ;
        RECT 2.37 0.71 2.49 1.17 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.465 ;
        RECT 1.875 1.31 2.25 1.445 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 0.76 0.585 1 ;
        RECT 0.305 0.83 0.565 1.09 ;
    END
  END A0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.61 1.265 2.85 1.385 ;
        RECT 2.68 0.885 2.83 1.145 ;
        RECT 2.68 0.885 2.8 1.385 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 0.825 1.725 1.09 ;
        RECT 1.45 0.76 1.69 1.005 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3384 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.885 3.12 1.145 ;
        RECT 2.515 1.505 3.09 1.625 ;
        RECT 2.97 0.47 3.09 1.625 ;
        RECT 2.85 0.4 2.97 0.64 ;
        RECT 1.255 0.47 3.09 0.59 ;
        RECT 2.515 1.505 2.635 1.865 ;
        RECT 1.255 0.4 1.375 0.64 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 1.99 -0.18 2.23 0.35 ;
        RECT 0.285 -0.18 0.405 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 0.985 2.135 1.105 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.055 1.985 2.875 1.985 2.875 2.105 1.315 2.105 1.315 1.925 1.195 1.925 1.195 1.805 1.435 1.805 1.435 1.985 2.095 1.985 2.095 1.745 2.215 1.745 2.215 1.985 2.755 1.985 2.755 1.865 2.935 1.865 2.935 1.745 3.055 1.745 ;
      POLYGON 1.795 1.865 1.675 1.865 1.675 1.685 0.625 1.685 0.625 1.83 0.505 1.83 0.505 1.565 1.795 1.565 ;
  END
END AOI222XL

MACRO OR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X6 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.95 2.135 1.13 ;
        RECT 1.755 0.94 2.015 1.13 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.25 2.595 1.37 ;
        RECT 2.475 0.94 2.595 1.37 ;
        RECT 2.335 0.94 2.595 1.09 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.49 2.955 1.61 ;
        RECT 2.835 1.105 2.955 1.61 ;
        RECT 0.68 1.28 1.075 1.61 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.155 1.465 3.41 1.725 ;
        RECT 0.41 1.73 3.38 1.85 ;
        RECT 3.155 1.465 3.38 1.85 ;
        RECT 3.155 1.22 3.275 1.85 ;
        RECT 0.41 1.22 0.53 1.85 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.735 0.4 5.855 0.915 ;
        RECT 5.555 0.795 5.855 0.915 ;
        RECT 3.995 0.91 5.675 1.03 ;
        RECT 5.535 1.39 5.655 2.21 ;
        RECT 3.855 1.39 5.655 1.51 ;
        RECT 4.935 1.175 5.15 1.51 ;
        RECT 4.935 0.91 5.055 1.51 ;
        RECT 4.895 0.4 5.015 1.03 ;
        RECT 4.695 1.39 4.815 2.21 ;
        RECT 3.995 0.4 4.115 1.03 ;
        RECT 3.855 1.39 3.975 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.315 -0.18 5.435 0.79 ;
        RECT 4.475 -0.18 4.595 0.79 ;
        RECT 3.515 0.46 3.755 0.58 ;
        RECT 3.515 -0.18 3.635 0.58 ;
        RECT 2.675 0.46 2.915 0.58 ;
        RECT 2.675 -0.18 2.795 0.58 ;
        RECT 1.835 0.46 2.075 0.58 ;
        RECT 1.835 -0.18 1.955 0.58 ;
        RECT 0.995 0.46 1.235 0.58 ;
        RECT 0.995 -0.18 1.115 0.58 ;
        RECT 0.215 -0.18 0.335 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.115 1.63 5.235 2.79 ;
        RECT 4.275 1.63 4.395 2.79 ;
        RECT 3.315 2.21 3.555 2.79 ;
        RECT 0.415 1.97 0.535 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.815 1.27 3.65 1.27 3.65 2.09 2.175 2.09 2.175 2.15 1.935 2.15 1.935 1.97 3.53 1.97 3.53 0.82 0.695 0.82 0.695 0.77 0.575 0.77 0.575 0.65 0.815 0.65 0.815 0.7 1.415 0.7 1.415 0.65 1.655 0.65 1.655 0.7 2.255 0.7 2.255 0.65 2.495 0.65 2.495 0.7 3.095 0.7 3.095 0.65 3.335 0.65 3.335 0.7 3.65 0.7 3.65 1.15 4.815 1.15 ;
  END
END OR4X6

MACRO ACHCONX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ACHCONX2 0 0 ;
  SIZE 14.5 BY 2.61 ;
  SYMMETRY X Y R90 ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.194 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.54 1.08 14.06 1.32 ;
        RECT 13.645 1.08 13.905 1.38 ;
    END
  END CI
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7841 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.72 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.089 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.165 1.13 3.51 1.49 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.194 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 1.23 0.565 1.38 ;
        RECT 0.19 0.975 0.43 1.38 ;
    END
  END A
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1716 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.97 1.57 12.93 1.69 ;
        RECT 10.53 0.36 12.93 0.48 ;
        RECT 11.905 1.23 12.165 1.38 ;
        RECT 10.53 1.805 12.09 1.925 ;
        RECT 11.97 0.36 12.09 1.925 ;
    END
  END CON
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.5 2.79 ;
        RECT 14.16 1.71 14.4 2.79 ;
        RECT 13.08 2.14 13.32 2.79 ;
        RECT 10.14 2.29 10.38 2.79 ;
        RECT 9.06 2.29 9.3 2.79 ;
        RECT 3.33 2.29 3.57 2.79 ;
        RECT 2.25 2.29 2.49 2.79 ;
        RECT 1.17 1.71 1.41 2.79 ;
        RECT 0.09 1.77 0.33 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.5 0.18 ;
        RECT 14.16 -0.18 14.4 0.725 ;
        RECT 13.08 -0.18 13.32 0.58 ;
        RECT 10.14 -0.18 10.38 0.32 ;
        RECT 9.06 -0.18 9.3 0.32 ;
        RECT 3.33 -0.18 3.57 0.32 ;
        RECT 2.25 -0.18 2.49 0.32 ;
        RECT 1.17 -0.18 1.41 0.64 ;
        RECT 0.09 -0.18 0.33 0.64 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 13.86 0.56 13.74 0.56 13.74 0.86 13.17 0.86 13.17 1.655 13.86 1.655 13.86 2.15 13.62 2.15 13.62 1.775 13.17 1.775 13.17 1.93 12.39 1.93 12.39 2.25 12.15 2.25 12.15 2.13 12.21 2.13 12.21 1.81 13.05 1.81 13.05 0.86 12.39 0.86 12.39 0.92 12.21 0.92 12.21 0.68 12.39 0.68 12.39 0.74 13.62 0.74 13.62 0.44 13.86 0.44 ;
      POLYGON 11.85 1.095 11.66 1.095 11.66 1.33 11 1.33 11 1.41 10.88 1.41 10.88 1.685 10.41 1.685 10.41 1.93 9.33 1.93 9.33 1.77 6.48 1.77 6.48 1.53 5.34 1.53 5.34 1.41 5.43 1.41 5.43 0.72 5.34 0.72 5.34 0.6 7.05 0.6 7.05 0.72 5.55 0.72 5.55 1.41 6.6 1.41 6.6 1.65 9.45 1.65 9.45 1.81 10.29 1.81 10.29 1.565 10.76 1.565 10.76 1.21 11.54 1.21 11.54 0.785 11.85 0.785 ;
      POLYGON 11.31 0.72 10.64 0.72 10.64 1.28 9.84 1.28 9.84 1.69 9.6 1.69 9.6 1.57 9.72 1.57 9.72 0.86 9.6 0.86 9.6 0.74 9.84 0.74 9.84 1.16 10.52 1.16 10.52 0.6 11.31 0.6 ;
      POLYGON 11.31 2.17 9.84 2.17 9.84 2.25 9.6 2.25 9.6 2.05 11.31 2.05 ;
      POLYGON 10.4 0.985 10.16 0.985 10.16 0.56 9.48 0.56 9.48 0.72 8.31 0.72 8.31 1.41 8.37 1.41 8.37 1.53 8.13 1.53 8.13 1.41 8.19 1.41 8.19 0.72 8.13 0.72 8.13 0.6 9.36 0.6 9.36 0.44 10.28 0.44 10.28 0.865 10.4 0.865 ;
      POLYGON 9.415 1.425 8.875 1.425 8.875 0.985 8.655 0.985 8.655 0.865 8.995 0.865 8.995 1.305 9.165 1.305 9.165 0.985 9.415 0.985 ;
      POLYGON 8.91 0.48 8.01 0.48 8.01 1.53 7.37 1.53 7.37 1.41 7.89 1.41 7.89 0.48 6.27 0.48 6.27 0.36 8.91 0.36 ;
      POLYGON 8.91 2.25 3.69 2.25 3.69 2.17 2.135 2.17 2.135 2.25 1.71 2.25 1.71 2.13 1.77 2.13 1.77 0.685 1.71 0.685 1.71 0.565 1.95 0.565 1.95 0.685 1.89 0.685 1.89 2.13 2.015 2.13 2.015 2.05 3.81 2.05 3.81 2.13 8.91 2.13 ;
      POLYGON 8.37 2.01 6.24 2.01 6.24 1.77 4.165 1.77 4.165 1.685 4 1.685 4 1.05 4.08 1.05 4.08 0.6 4.5 0.6 4.5 0.72 4.2 0.72 4.2 1.17 4.12 1.17 4.12 1.565 4.285 1.565 4.285 1.65 6.36 1.65 6.36 1.89 8.37 1.89 ;
      POLYGON 7.77 1.29 7.55 1.29 7.55 1.125 6.98 1.125 6.98 0.96 6.325 0.96 6.325 0.84 7.1 0.84 7.1 1.005 7.77 1.005 ;
      POLYGON 7.03 1.49 6.79 1.49 6.79 1.365 6.715 1.365 6.715 1.29 5.8 1.29 5.8 1.025 5.68 1.025 5.68 0.84 5.92 0.84 5.92 1.17 6.835 1.17 6.835 1.245 7.03 1.245 ;
      POLYGON 6.12 0.48 3.96 0.48 3.96 0.56 2.385 0.56 2.385 1.81 4.045 1.81 4.045 1.89 6.12 1.89 6.12 2.01 3.925 2.01 3.925 1.93 2.265 1.93 2.265 1.25 2.05 1.25 2.05 1.13 2.265 1.13 2.265 0.44 3.72 0.44 3.72 0.36 6.12 0.36 ;
      POLYGON 5.08 1.425 4.24 1.425 4.24 1.305 4.96 1.305 4.96 1.025 4.9 1.025 4.9 0.73 5.08 0.73 ;
      POLYGON 3.88 0.985 3.64 0.985 3.64 0.875 2.97 0.875 2.97 1.57 3.03 1.57 3.03 1.69 2.79 1.69 2.79 1.57 2.85 1.57 2.85 0.875 2.79 0.875 2.79 0.74 3.03 0.74 3.03 0.755 3.88 0.755 ;
      POLYGON 1.51 1.25 0.81 1.25 0.81 1.625 0.87 1.625 0.87 2.065 0.63 2.065 0.63 1.625 0.69 1.625 0.69 0.685 0.63 0.685 0.63 0.565 0.87 0.565 0.87 0.685 0.81 0.685 0.81 1.13 1.51 1.13 ;
  END
END ACHCONX2

MACRO XOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3XL 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3684 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.27 1.56 8.51 2.25 ;
        RECT 8.39 0.36 8.51 2.25 ;
        RECT 8.135 0.65 8.51 0.8 ;
        RECT 8.27 0.36 8.51 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.084 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.07 0.325 1.47 ;
        RECT 0.07 1.175 0.325 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3168 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.2571 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.23 1.145 1.38 ;
        RECT 0.845 1.03 1.025 1.375 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 1.35 6.81 1.47 ;
        RECT 6.08 1.23 6.365 1.47 ;
        RECT 6.08 0.905 6.2 1.47 ;
        RECT 5.695 0.905 6.2 1.025 ;
    END
  END C
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.73 2.29 7.97 2.79 ;
        RECT 7.79 1.69 7.91 2.79 ;
        RECT 1.865 2.27 2.105 2.79 ;
        RECT 0.685 2.29 0.925 2.79 ;
        RECT 0.745 1.97 0.865 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.73 -0.18 7.97 0.32 ;
        RECT 7.79 -0.18 7.91 0.67 ;
        RECT 1.865 -0.18 2.105 0.32 ;
        RECT 0.685 -0.18 0.925 0.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.23 1.315 7.67 1.315 7.67 2.17 6.26 2.17 6.26 1.89 6.56 1.89 6.56 2.05 7.55 2.05 7.55 0.62 7.42 0.62 7.42 0.48 6.26 0.48 6.26 0.36 7.54 0.36 7.54 0.5 7.67 0.5 7.67 1.195 7.99 1.195 7.99 1.075 8.23 1.075 ;
      POLYGON 7.43 0.86 7.345 0.86 7.345 1.81 7.43 1.81 7.43 1.93 7.19 1.93 7.19 1.81 7.225 1.81 7.225 0.86 7.19 0.86 7.19 0.74 7.43 0.74 ;
      POLYGON 7.05 1.77 7.04 1.77 7.04 1.79 6.8 1.79 6.8 1.77 4.275 1.77 4.275 1.65 5.095 1.65 5.095 0.72 4.27 0.72 4.27 0.6 5.215 0.6 5.215 1.65 6.93 1.65 6.93 0.72 6.8 0.72 6.8 0.6 7.05 0.6 ;
      POLYGON 5.96 0.705 5.9 0.705 5.9 0.72 5.48 0.72 5.48 1.405 5.96 1.405 5.96 1.525 5.36 1.525 5.36 0.6 5.72 0.6 5.72 0.585 5.96 0.585 ;
      RECT 2.985 1.89 5.96 2.01 ;
      RECT 2.405 0.36 5.64 0.48 ;
      RECT 2.405 2.13 5.64 2.25 ;
      POLYGON 4.84 1.04 4.17 1.04 4.17 1.415 4.05 1.415 4.05 0.92 4.84 0.92 ;
      POLYGON 3.985 0.72 3.84 0.72 3.84 1.77 1.725 1.77 1.725 2.17 0.985 2.17 0.985 1.81 0.325 1.81 0.325 1.93 0.145 1.93 0.145 1.69 0.505 1.69 0.505 0.92 0.205 0.92 0.205 0.44 1.605 0.44 1.605 0.32 1.725 0.32 1.725 0.56 0.325 0.56 0.325 0.8 0.625 0.8 0.625 1.69 1.105 1.69 1.105 2.05 1.605 2.05 1.605 1.65 3.72 1.65 3.72 0.6 3.985 0.6 ;
      POLYGON 3.585 1.04 3.405 1.04 3.405 1 2.81 1 2.81 1.16 2.885 1.16 2.885 1.28 2.645 1.28 2.645 1.16 2.69 1.16 2.69 0.88 3.405 0.88 3.405 0.8 3.585 0.8 ;
      POLYGON 3.225 1.53 1.94 1.53 1.94 0.6 3.205 0.6 3.205 0.72 2.06 0.72 2.06 1.41 3.225 1.41 ;
      POLYGON 1.485 1.12 1.405 1.12 1.405 1.81 1.465 1.81 1.465 1.93 1.225 1.93 1.225 1.81 1.285 1.81 1.285 1.12 1.245 1.12 1.245 1 1.285 1 1.285 0.8 1.225 0.8 1.225 0.68 1.465 0.68 1.465 0.8 1.405 0.8 1.405 1 1.485 1 ;
  END
END XOR3XL

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.03 1.38 1.485 ;
        RECT 1.23 1 1.35 1.485 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.2 1.085 1.32 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1 0.51 1.485 ;
        RECT 0.36 1 0.51 1.455 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3284 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.065 1.605 1.67 1.725 ;
        RECT 1.5 1.465 1.67 1.725 ;
        RECT 1.5 0.71 1.62 1.725 ;
        RECT 1.485 0.59 1.605 0.83 ;
        RECT 1.065 1.605 1.185 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.645 -0.18 0.765 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.485 1.845 1.605 2.79 ;
        RECT 0.425 1.605 0.545 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.185 0.88 0.225 0.88 0.225 0.59 0.345 0.59 0.345 0.76 1.065 0.76 1.065 0.59 1.185 0.59 ;
  END
END OAI21X1

MACRO DLY3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.315 0.68 5.555 0.8 ;
        RECT 5.375 0.68 5.495 2.21 ;
        RECT 4.42 0.885 5.495 1.005 ;
        RECT 5.315 0.68 5.495 1.005 ;
        RECT 4.535 0.885 4.655 2.21 ;
        RECT 4.42 0.68 4.595 1.145 ;
        RECT 4.355 0.68 4.595 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.885 2.86 1.145 ;
        RECT 2.605 1.025 2.78 1.265 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.57 0.92 8.69 1.74 ;
        RECT 8.435 0.92 8.69 1.04 ;
        RECT 8.435 -0.18 8.555 1.04 ;
        RECT 7.735 0.6 7.975 0.72 ;
        RECT 7.835 -0.18 7.955 0.72 ;
        RECT 6.455 1.24 6.635 1.48 ;
        RECT 6.515 -0.18 6.635 1.48 ;
        RECT 5.915 0.68 6.155 0.8 ;
        RECT 5.915 -0.18 6.035 0.8 ;
        RECT 4.835 -0.18 5.075 0.32 ;
        RECT 3.875 -0.18 3.995 0.53 ;
        RECT 3.625 1.04 3.745 1.42 ;
        RECT 3.315 1.04 3.745 1.16 ;
        RECT 3.315 -0.18 3.435 1.16 ;
        RECT 2.595 -0.18 2.835 0.34 ;
        RECT 1.655 1.37 1.895 1.49 ;
        RECT 1.775 0.76 1.895 1.49 ;
        RECT 1.575 0.76 1.895 0.88 ;
        RECT 1.575 -0.18 1.695 0.88 ;
        RECT 1.175 -0.18 1.295 0.64 ;
        RECT 0.375 -0.18 0.495 1.36 ;
        RECT 0.355 1.24 0.475 1.48 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.33 1.16 8.45 1.4 ;
        RECT 7.37 1.16 8.45 1.28 ;
        RECT 7.37 1.76 7.61 2.79 ;
        RECT 7.37 1.08 7.49 2.79 ;
        RECT 7.235 1.08 7.49 1.2 ;
        RECT 5.795 1.58 5.915 2.79 ;
        RECT 4.955 1.56 5.075 2.79 ;
        RECT 4.115 1.93 4.235 2.79 ;
        RECT 3.225 1.28 3.465 1.4 ;
        RECT 3.225 1.28 3.345 2.79 ;
        RECT 2.785 1.66 2.905 2.79 ;
        RECT 0.615 1 1.655 1.12 ;
        RECT 1.175 1.61 1.535 1.73 ;
        RECT 1.415 1 1.535 1.73 ;
        RECT 0.975 1.84 1.295 2.79 ;
        RECT 1.175 1.61 1.295 2.79 ;
        RECT 0.855 1.84 1.295 1.96 ;
        RECT 0.615 0.78 0.855 1.12 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.93 2.02 8.41 2.02 8.41 1.98 8.33 1.98 8.33 1.64 7.69 1.64 7.69 1.4 7.93 1.4 7.93 1.52 8.45 1.52 8.45 1.86 8.81 1.86 8.81 0.8 8.675 0.8 8.675 0.68 8.93 0.68 ;
      POLYGON 8.315 0.48 8.215 0.48 8.215 0.96 7.495 0.96 7.495 0.62 6.875 0.62 6.875 1.72 6.555 1.72 6.555 1.84 6.435 1.84 6.435 1.6 6.755 1.6 6.755 0.5 7.615 0.5 7.615 0.84 8.095 0.84 8.095 0.48 8.075 0.48 8.075 0.36 8.315 0.36 ;
      POLYGON 7.375 0.86 7.255 0.86 7.255 0.96 7.115 0.96 7.115 1.56 7.19 1.56 7.19 2.21 7.07 2.21 7.07 2.08 6.035 2.08 6.035 1.42 5.615 1.42 5.615 1.3 6.155 1.3 6.155 1.96 6.995 1.96 6.995 0.84 7.135 0.84 7.135 0.74 7.375 0.74 ;
      POLYGON 6.395 1.04 5.675 1.04 5.675 0.56 4.235 0.56 4.235 0.77 3.985 0.77 3.985 1.66 3.905 1.66 3.905 1.78 3.785 1.78 3.785 1.54 3.865 1.54 3.865 0.92 3.555 0.92 3.555 0.65 4.115 0.65 4.115 0.44 5.795 0.44 5.795 0.92 6.275 0.92 6.275 0.48 6.155 0.48 6.155 0.36 6.395 0.36 ;
      POLYGON 3.195 0.54 3.075 0.54 3.075 0.58 2.135 0.58 2.135 1.73 2.095 1.73 2.095 1.87 1.975 1.87 1.975 1.61 2.015 1.61 2.015 0.64 1.815 0.64 1.815 0.4 1.935 0.4 1.935 0.46 2.955 0.46 2.955 0.42 3.195 0.42 ;
      POLYGON 2.495 0.86 2.485 0.86 2.485 2.11 1.655 2.11 1.655 2.25 1.415 2.25 1.415 2.13 1.535 2.13 1.535 1.99 2.365 1.99 2.365 0.86 2.255 0.86 2.255 0.74 2.495 0.74 ;
      POLYGON 1.295 1.49 1.055 1.49 1.055 1.72 0.395 1.72 0.395 1.81 0.115 1.81 0.115 0.52 0.135 0.52 0.135 0.4 0.255 0.4 0.255 0.64 0.235 0.64 0.235 1.6 0.935 1.6 0.935 1.37 1.295 1.37 ;
  END
END DLY3X4

MACRO TLATNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX2 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.615 1.16 0.835 1.51 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.33 3.12 1.725 ;
        RECT 2.88 1.33 3.12 1.45 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.69 1.09 4.86 1.5 ;
        RECT 4.69 1.09 4.81 1.515 ;
    END
  END SN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.67 1 7.81 1.27 ;
        RECT 7.61 0.86 7.78 1.145 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.33 0.68 5.45 1.025 ;
        RECT 5.27 1.38 5.39 1.67 ;
        RECT 5.32 0.885 5.44 1.5 ;
        RECT 5.29 0.885 5.44 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.19 1.145 7.31 1.67 ;
        RECT 7.06 1.145 7.31 1.265 ;
        RECT 7.03 0.885 7.18 1.145 ;
        RECT 7.01 0.68 7.13 1.025 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.43 -0.18 7.55 0.73 ;
        RECT 6.59 -0.18 6.71 0.73 ;
        RECT 5.75 -0.18 5.87 0.73 ;
        RECT 4.91 -0.18 5.03 0.73 ;
        RECT 2.715 0.61 2.955 0.73 ;
        RECT 2.715 -0.18 2.835 0.73 ;
        RECT 0.495 0.68 0.735 0.8 ;
        RECT 0.495 -0.18 0.615 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.67 2.03 7.79 2.79 ;
        RECT 6.65 2.03 6.89 2.15 ;
        RECT 6.65 2.03 6.77 2.79 ;
        RECT 5.69 2.03 5.93 2.15 ;
        RECT 5.69 2.03 5.81 2.79 ;
        RECT 4.79 2.23 4.91 2.79 ;
        RECT 4.29 2.23 4.41 2.79 ;
        RECT 3.15 2.23 3.27 2.79 ;
        RECT 2.245 2.29 2.485 2.79 ;
        RECT 0.615 1.87 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.27 1.79 7.88 1.79 7.88 1.91 5.495 1.91 5.495 2.11 4.17 2.11 4.17 2.25 3.61 2.25 3.61 2.13 4.05 2.13 4.05 1.99 5.375 1.99 5.375 1.79 7.76 1.79 7.76 1.67 8.15 1.67 8.15 1.55 7.93 1.55 7.93 0.68 8.05 0.68 8.05 1.43 8.27 1.43 ;
      POLYGON 6.91 1.29 6.35 1.29 6.35 1.67 6.23 1.67 6.23 0.92 6.17 0.92 6.17 0.68 6.29 0.68 6.29 0.8 6.35 0.8 6.35 1.17 6.91 1.17 ;
      POLYGON 5.17 1.26 5.05 1.26 5.05 0.97 4.55 0.97 4.55 1.87 4.43 1.87 4.43 0.97 4.21 0.97 4.21 0.58 3.945 0.58 3.945 0.5 3.27 0.5 3.27 0.97 2.275 0.97 2.275 0.48 2.155 0.48 2.155 0.36 2.395 0.36 2.395 0.85 3.15 0.85 3.15 0.38 4.065 0.38 4.065 0.46 4.33 0.46 4.33 0.85 5.17 0.85 ;
      POLYGON 4.27 1.87 3.93 1.87 3.93 2.01 3.205 2.01 3.205 2.11 2.94 2.11 2.94 2.17 1.495 2.17 1.495 1.75 1.615 1.75 1.615 1.57 1.655 1.57 1.655 0.62 1.775 0.62 1.775 1.69 1.735 1.69 1.735 1.87 1.615 1.87 1.615 2.05 2.82 2.05 2.82 1.99 3.085 1.99 3.085 1.89 3.81 1.89 3.81 1.75 4.15 1.75 4.15 1.11 4.27 1.11 ;
      POLYGON 3.69 1.77 3.45 1.77 3.45 1.21 1.915 1.21 1.915 0.5 1.535 0.5 1.535 1.45 1.415 1.45 1.415 1.04 0.495 1.04 0.495 1.22 0.355 1.22 0.355 0.98 0.375 0.98 0.375 0.92 1.415 0.92 1.415 0.38 2.035 0.38 2.035 1.02 2.155 1.02 2.155 1.09 3.475 1.09 3.475 0.62 3.595 0.62 3.595 1.21 3.57 1.21 3.57 1.65 3.69 1.65 ;
      POLYGON 2.85 1.87 2.095 1.87 2.095 1.93 1.855 1.93 1.855 1.81 1.975 1.81 1.975 1.75 2.85 1.75 ;
      POLYGON 1.235 1.28 1.075 1.28 1.075 1.75 0.315 1.75 0.315 1.99 0.195 1.99 0.195 1.87 0.115 1.87 0.115 0.74 0.135 0.74 0.135 0.62 0.255 0.62 0.255 0.86 0.235 0.86 0.235 1.63 0.955 1.63 0.955 1.16 1.235 1.16 ;
  END
END TLATNSRX2

MACRO AND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.04 0.51 1.5 ;
        RECT 0.36 1.04 0.48 1.53 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 1.04 0.89 1.35 ;
        RECT 0.65 1.12 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.25 1.465 1.67 1.585 ;
        RECT 1.25 1.345 1.37 1.585 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.175 1.96 1.435 ;
        RECT 1.83 1.175 1.95 2.01 ;
        RECT 1.81 0.68 1.93 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.39 -0.18 1.51 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.41 1.89 1.53 2.79 ;
        RECT 0.57 1.89 0.69 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 1.34 1.57 1.34 1.57 1.225 1.13 1.225 1.13 1.825 1.11 1.825 1.11 2.01 0.99 2.01 0.99 1.77 0.33 1.77 0.33 1.95 0.09 1.95 0.09 1.83 0.21 1.83 0.21 1.65 1.01 1.65 1.01 0.92 0.29 0.92 0.29 0.68 0.41 0.68 0.41 0.8 1.13 0.8 1.13 1.105 1.57 1.105 1.57 1.1 1.69 1.1 ;
  END
END AND3XL

MACRO DFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSXL 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.135 1.22 3.465 1.435 ;
        RECT 3.015 1.22 3.465 1.41 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.035 1.22 8.155 1.51 ;
        RECT 7.9 1.175 8.05 1.475 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 1.04 8.63 1.435 ;
        RECT 8.48 0.835 8.6 1.435 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.66 1.485 1.58 ;
        RECT 1.23 0.885 1.485 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.375 -0.18 8.495 0.38 ;
        RECT 6.605 -0.18 6.845 0.32 ;
        RECT 3.295 -0.18 3.415 0.4 ;
        RECT 1.845 -0.18 1.965 0.38 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.195 1.68 8.315 2.79 ;
        RECT 6.955 2.2 7.075 2.79 ;
        RECT 4.375 2.29 4.615 2.79 ;
        RECT 3.475 2.05 3.595 2.79 ;
        RECT 2.515 1.73 2.635 2.79 ;
        RECT 1.845 1.98 1.965 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.87 1.675 8.735 1.675 8.735 1.8 8.615 1.8 8.615 1.555 8.75 1.555 8.75 0.9 8.735 0.9 8.735 0.66 8.135 0.66 8.135 0.54 7.515 0.54 7.515 1.46 7.395 1.46 7.395 0.56 5.675 0.56 5.675 1.46 5.555 1.46 5.555 0.56 5.195 0.56 5.195 0.52 5.075 0.52 5.075 0.4 5.315 0.4 5.315 0.44 6.245 0.44 6.245 0.4 6.485 0.4 6.485 0.44 7.395 0.44 7.395 0.42 7.755 0.42 7.755 0.4 7.995 0.4 7.995 0.42 8.255 0.42 8.255 0.54 8.855 0.54 8.855 0.78 8.87 0.78 ;
      POLYGON 7.755 1.7 7.675 1.7 7.675 1.94 6.835 1.94 6.835 2.22 4.735 2.22 4.735 2.17 4.055 2.17 4.055 2.05 4.855 2.05 4.855 2.1 6.715 2.1 6.715 1.82 7.555 1.82 7.555 1.58 7.635 1.58 7.635 0.66 7.755 0.66 ;
      POLYGON 7.195 1.46 7.075 1.46 7.075 1.18 6.245 1.18 6.245 1.62 6.355 1.62 6.355 1.74 6.115 1.74 6.115 1.62 6.125 1.62 6.125 1.26 6.035 1.26 6.035 1.02 6.125 1.02 6.125 0.72 6.365 0.72 6.365 0.84 6.245 0.84 6.245 1.06 7.195 1.06 ;
      POLYGON 6.915 1.42 6.795 1.42 6.795 1.7 6.595 1.7 6.595 1.98 5.785 1.98 5.785 1.96 5.065 1.96 5.065 1.6 4.8 1.6 4.8 1.57 4.135 1.57 4.135 1.69 3.895 1.69 3.895 1.57 4.015 1.57 4.015 1.45 4.275 1.45 4.275 0.68 4.395 0.68 4.395 1.45 4.92 1.45 4.92 1.48 5.185 1.48 5.185 1.84 5.785 1.84 5.785 1.58 5.795 1.58 5.795 0.68 5.915 0.68 5.915 1.7 5.905 1.7 5.905 1.86 6.475 1.86 6.475 1.58 6.675 1.58 6.675 1.3 6.915 1.3 ;
      POLYGON 5.545 1.72 5.305 1.72 5.305 1.16 4.515 1.16 4.515 0.56 4.155 0.56 4.155 0.72 4.035 0.72 4.035 1.1 2.185 1.1 2.185 1.22 2.065 1.22 2.065 0.98 3.915 0.98 3.915 0.6 4.035 0.6 4.035 0.44 4.635 0.44 4.635 1.04 5.305 1.04 5.305 0.86 5.195 0.86 5.195 0.74 5.435 0.74 5.435 0.86 5.425 0.86 5.425 1.6 5.545 1.6 ;
      POLYGON 4.955 0.92 4.835 0.92 4.835 0.72 4.755 0.72 4.755 0.36 4.875 0.36 4.875 0.6 4.955 0.6 ;
      POLYGON 4.945 1.84 4.825 1.84 4.825 1.93 2.995 1.93 2.995 1.63 3.115 1.63 3.115 1.81 4.705 1.81 4.705 1.72 4.945 1.72 ;
      POLYGON 3.915 0.48 3.795 0.48 3.795 0.74 2.775 0.74 2.775 0.86 2.535 0.86 2.535 0.74 2.655 0.74 2.655 0.62 3.675 0.62 3.675 0.36 3.915 0.36 ;
      POLYGON 2.895 1.37 2.425 1.37 2.425 1.46 2.325 1.46 2.325 1.58 2.205 1.58 2.205 1.46 1.825 1.46 1.825 1.2 1.605 1.2 1.605 1.08 1.825 1.08 1.825 0.72 2.385 0.72 2.385 0.84 1.945 0.84 1.945 1.34 2.305 1.34 2.305 1.25 2.895 1.25 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END DFFSXL

MACRO NAND4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBXL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.94 0.395 1.18 ;
        RECT 0.07 0.94 0.395 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.425 1.32 2.665 1.505 ;
        RECT 2.335 1.23 2.595 1.44 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.52 ;
        RECT 1.425 1.325 1.545 1.67 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.23 1.145 1.5 ;
        RECT 0.815 1.36 1.055 1.61 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2976 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.945 0.695 2.065 2.09 ;
        RECT 1.105 1.79 2.065 1.91 ;
        RECT 1.81 1.465 2.065 1.91 ;
        RECT 1.005 0.695 2.065 0.815 ;
        RECT 1.105 1.79 1.225 2.09 ;
        RECT 0.885 0.595 1.125 0.715 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.325 -0.18 2.445 0.775 ;
        RECT 0.135 -0.18 0.255 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.365 1.97 2.485 2.79 ;
        RECT 1.465 2.03 1.705 2.15 ;
        RECT 1.465 2.03 1.585 2.79 ;
        RECT 0.685 1.97 0.805 2.79 ;
        RECT 0.135 1.46 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.925 0.715 2.905 0.715 2.905 2.09 2.785 2.09 2.785 1.11 2.185 1.11 2.185 0.99 2.785 0.99 2.785 0.715 2.685 0.715 2.685 0.595 2.925 0.595 ;
      POLYGON 1.825 1.055 0.675 1.055 0.675 1.58 0.555 1.58 0.555 0.525 0.675 0.525 0.675 0.935 1.825 0.935 ;
  END
END NAND4BBXL

MACRO CLKBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX16 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.685 1.26 7.285 1.38 ;
        RECT 6.685 1.23 6.945 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.565 0.715 5.805 0.835 ;
        RECT 5.625 1.295 5.745 2.21 ;
        RECT 0.545 0.765 5.685 0.885 ;
        RECT 0.545 1.295 5.745 1.415 ;
        RECT 4.725 0.715 4.965 0.885 ;
        RECT 4.785 1.295 4.905 2.21 ;
        RECT 3.885 0.715 4.125 0.885 ;
        RECT 3.945 1.295 4.065 2.21 ;
        RECT 3.045 0.715 3.285 0.885 ;
        RECT 3.105 1.295 3.225 2.21 ;
        RECT 2.205 0.715 2.445 0.885 ;
        RECT 2.265 1.295 2.385 2.21 ;
        RECT 1.365 0.715 1.605 0.885 ;
        RECT 1.425 1.295 1.545 2.21 ;
        RECT 0.585 1.295 0.8 1.725 ;
        RECT 0.585 1.295 0.705 2.21 ;
        RECT 0.585 0.645 0.705 0.885 ;
        RECT 0.545 0.765 0.665 1.415 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.725 -0.18 7.845 0.705 ;
        RECT 6.885 -0.18 7.005 0.705 ;
        RECT 6.045 -0.18 6.165 0.705 ;
        RECT 5.205 -0.18 5.325 0.645 ;
        RECT 4.365 -0.18 4.485 0.645 ;
        RECT 3.525 -0.18 3.645 0.645 ;
        RECT 2.685 -0.18 2.805 0.645 ;
        RECT 1.845 -0.18 1.965 0.645 ;
        RECT 1.005 -0.18 1.125 0.64 ;
        RECT 0.165 -0.18 0.285 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.725 1.56 7.845 2.79 ;
        RECT 6.885 1.74 7.005 2.79 ;
        RECT 6.045 1.56 6.165 2.79 ;
        RECT 5.205 1.535 5.325 2.79 ;
        RECT 4.365 1.535 4.485 2.79 ;
        RECT 3.525 1.535 3.645 2.79 ;
        RECT 2.685 1.535 2.805 2.79 ;
        RECT 1.845 1.535 1.965 2.79 ;
        RECT 1.005 1.535 1.125 2.79 ;
        RECT 0.165 1.465 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.425 0.945 6.565 0.945 6.565 1.5 7.425 1.5 7.425 2.21 7.305 2.21 7.305 1.62 6.585 1.62 6.585 2.21 6.465 2.21 6.465 1.62 6.445 1.62 6.445 1.175 0.785 1.175 0.785 1.055 6.445 1.055 6.445 0.825 6.465 0.825 6.465 0.655 6.585 0.655 6.585 0.825 7.305 0.825 7.305 0.655 7.425 0.655 ;
  END
END CLKBUFX16

MACRO OAI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X1 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.985 2.54 1.44 ;
        RECT 2.405 0.895 2.525 1.44 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 1 2.005 1.35 ;
        RECT 1.81 1.085 1.96 1.435 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.14 1.09 1.435 ;
        RECT 0.835 1.1 0.955 1.38 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.035 1.67 1.49 ;
        RECT 1.545 1.01 1.665 1.49 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.01 0.51 1.495 ;
        RECT 0.36 1.01 0.51 1.465 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7639 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.385 1.61 2.78 1.73 ;
        RECT 2.66 0.745 2.78 1.73 ;
        RECT 2.645 0.6 2.765 0.865 ;
        RECT 2.445 1.56 2.78 1.73 ;
        RECT 2.445 1.56 2.565 2.21 ;
        RECT 2.39 1.61 2.565 2.015 ;
        RECT 1.385 1.61 1.505 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 0.995 -0.18 1.115 0.65 ;
        RECT 0.155 -0.18 0.275 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.025 1.85 2.145 2.79 ;
        RECT 0.355 1.615 0.475 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.345 0.65 2.225 0.65 2.225 0.53 2.045 0.53 2.045 0.48 1.505 0.48 1.505 0.65 1.385 0.65 1.385 0.36 2.165 0.36 2.165 0.41 2.345 0.41 ;
      POLYGON 1.925 0.88 1.765 0.88 1.765 0.89 0.575 0.89 0.575 0.6 0.695 0.6 0.695 0.77 1.645 0.77 1.645 0.76 1.805 0.76 1.805 0.6 1.925 0.6 ;
  END
END OAI221X1

MACRO AND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4XL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.23 0.565 1.5 ;
        RECT 0.325 1.1 0.565 1.5 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.095 1.09 1.46 ;
        RECT 0.815 1.095 0.935 1.465 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 1.095 1.38 1.56 ;
        RECT 1.21 1.095 1.33 1.59 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.37 1.96 1.725 ;
        RECT 1.74 1.215 1.86 1.575 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.355 0.855 2.475 1.83 ;
        RECT 2.13 0.855 2.475 0.975 ;
        RECT 2.1 0.595 2.25 0.855 ;
        RECT 1.935 0.595 2.25 0.735 ;
        RECT 1.935 0.495 2.055 0.735 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.515 -0.18 1.635 0.735 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.875 2.23 1.995 2.79 ;
        RECT 0.915 2.23 1.035 2.79 ;
        RECT 0.135 1.71 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.98 1.095 1.86 1.095 1.86 0.975 1.62 0.975 1.62 1.83 1.515 1.83 1.515 1.95 1.395 1.95 1.395 1.83 0.495 1.83 0.495 1.71 1.5 1.71 1.5 0.975 0.395 0.975 0.395 0.675 0.275 0.675 0.275 0.555 0.515 0.555 0.515 0.855 1.98 0.855 ;
  END
END AND4XL

MACRO OAI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.03 1.38 1.485 ;
        RECT 1.23 1 1.35 1.485 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.03 1.67 1.485 ;
        RECT 1.55 1 1.67 1.485 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.985 0.44 1.245 ;
        RECT 0.32 0.76 0.44 1.245 ;
        RECT 0.07 0.985 0.22 1.44 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.065 1.09 1.435 ;
        RECT 0.84 1.01 0.96 1.385 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3284 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.32 1.605 1.96 1.725 ;
        RECT 1.84 0.59 1.96 1.725 ;
        RECT 1.81 0.885 1.96 1.145 ;
        RECT 1.32 1.605 1.44 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1 -0.18 1.12 0.64 ;
        RECT 0.16 -0.18 0.28 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.74 1.845 1.86 2.79 ;
        RECT 0.36 1.56 0.48 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.54 0.88 0.58 0.88 0.58 0.59 0.7 0.59 0.7 0.76 1.42 0.76 1.42 0.59 1.54 0.59 ;
  END
END OAI31X1

MACRO OA21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.77 1.38 1.145 ;
        RECT 1.23 0.77 1.35 1.26 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.95 1.295 ;
        RECT 0.83 1.055 0.95 1.295 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.125 0.51 1.56 ;
        RECT 0.39 1.08 0.51 1.56 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 0.65 2.43 0.77 ;
        RECT 1.97 1.005 2.25 1.145 ;
        RECT 2.13 0.65 2.25 1.145 ;
        RECT 2.1 0.885 2.25 1.145 ;
        RECT 1.97 1.005 2.09 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.77 -0.18 1.89 0.53 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.55 1.62 1.67 2.79 ;
        RECT 0.35 1.68 0.47 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 1.48 1.62 1.48 1.62 1.5 1.19 1.5 1.19 1.8 1.07 1.8 1.07 1.38 1.5 1.38 1.5 0.68 1.62 0.68 1.62 1.24 1.82 1.24 ;
      POLYGON 1.11 0.92 0.99 0.92 0.99 0.86 0.075 0.86 0.075 0.74 0.99 0.74 0.99 0.68 1.11 0.68 ;
  END
END OA21X1

MACRO DLY4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X4 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 1.4 2.235 1.52 ;
        RECT 2.055 0.59 2.175 1.52 ;
        RECT 1.23 1.025 2.175 1.145 ;
        RECT 1.215 0.885 1.38 1.025 ;
        RECT 1.035 1.4 1.35 1.52 ;
        RECT 1.23 0.885 1.35 1.52 ;
        RECT 1.215 0.59 1.335 1.025 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.25 10.575 1.49 ;
        RECT 10.25 1.37 10.575 1.49 ;
        RECT 10.22 1.465 10.37 1.725 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.235 -0.18 10.355 0.89 ;
        RECT 9.685 1.24 9.955 1.36 ;
        RECT 9.835 -0.18 9.955 1.36 ;
        RECT 9.685 1.24 9.805 1.48 ;
        RECT 8.365 -0.18 8.485 0.38 ;
        RECT 7.585 -0.18 7.705 1.36 ;
        RECT 7.485 1.24 7.605 1.48 ;
        RECT 6.635 1.2 6.875 1.32 ;
        RECT 6.715 -0.18 6.835 1.32 ;
        RECT 6.015 -0.18 6.135 0.84 ;
        RECT 5.155 1.51 5.415 1.63 ;
        RECT 5.155 -0.18 5.275 1.63 ;
        RECT 4.135 1.48 4.555 1.72 ;
        RECT 4.435 0.98 4.555 1.72 ;
        RECT 4.225 0.98 4.555 1.1 ;
        RECT 4.225 -0.18 4.345 1.1 ;
        RECT 3.885 -0.18 4.005 0.86 ;
        RECT 3.075 1 3.195 1.24 ;
        RECT 2.815 1 3.195 1.12 ;
        RECT 2.815 -0.18 2.935 1.12 ;
        RECT 2.475 -0.18 2.595 0.64 ;
        RECT 1.635 -0.18 1.755 0.64 ;
        RECT 0.795 -0.18 0.915 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.245 2.23 10.365 2.79 ;
        RECT 8.945 1 9.065 1.24 ;
        RECT 7.825 1 9.065 1.12 ;
        RECT 8.425 1.68 8.545 2.79 ;
        RECT 7.965 1 8.085 2.79 ;
        RECT 7.825 1 8.085 1.24 ;
        RECT 6.195 2.16 6.315 2.79 ;
        RECT 6.075 2.16 6.315 2.28 ;
        RECT 4.995 1.79 5.115 2.79 ;
        RECT 3.515 2.08 3.755 2.2 ;
        RECT 3.515 2.08 3.635 2.79 ;
        RECT 2.535 1.88 2.655 2.79 ;
        RECT 1.515 1.88 1.755 2 ;
        RECT 1.515 1.88 1.635 2.79 ;
        RECT 0.555 1.88 0.795 2 ;
        RECT 0.555 1.88 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.845 1.85 10.725 1.85 10.725 1.73 10.695 1.73 10.695 1.13 10.335 1.13 10.335 1.17 10.075 1.17 10.075 1.05 10.215 1.05 10.215 1.01 10.655 1.01 10.655 0.65 10.775 0.65 10.775 0.89 10.815 0.89 10.815 1.61 10.845 1.61 ;
      POLYGON 9.715 0.89 9.565 0.89 9.565 1.6 9.665 1.6 9.665 1.84 9.545 1.84 9.545 1.72 9.445 1.72 9.445 0.77 9.595 0.77 9.595 0.65 9.56 0.65 9.56 0.54 8.765 0.54 8.765 0.52 8.645 0.52 8.645 0.4 8.885 0.4 8.885 0.42 9.68 0.42 9.68 0.53 9.715 0.53 ;
      POLYGON 9.325 1.48 9.185 1.48 9.185 1.8 9.065 1.8 9.065 1.48 8.205 1.48 8.205 1.24 8.325 1.24 8.325 1.36 9.205 1.36 9.205 0.66 9.325 0.66 ;
      POLYGON 7.845 1.8 6.055 1.8 6.055 1.77 6.015 1.77 6.015 1.53 6.055 1.53 6.055 0.96 6.295 0.96 6.295 0.36 6.535 0.36 6.535 1.08 6.175 1.08 6.175 1.68 7.245 1.68 7.245 0.78 7.345 0.78 7.345 0.66 7.465 0.66 7.465 0.9 7.365 0.9 7.365 1.68 7.845 1.68 ;
      POLYGON 7.115 1.56 6.295 1.56 6.295 1.44 6.995 1.44 6.995 1.08 6.955 1.08 6.955 0.62 7.075 0.62 7.075 0.96 7.115 0.96 ;
      POLYGON 7.015 2.04 5.775 2.04 5.775 0.48 5.395 0.48 5.395 0.36 5.895 0.36 5.895 1.92 7.015 1.92 ;
      POLYGON 5.655 1.87 5.555 1.87 5.555 2.09 5.435 2.09 5.435 1.75 5.535 1.75 5.535 1.13 5.655 1.13 ;
      POLYGON 5.035 0.86 4.915 0.86 4.915 0.48 4.775 0.48 4.775 0.36 5.035 0.36 ;
      POLYGON 4.795 1.97 4.395 1.97 4.395 2.09 4.275 2.09 4.275 1.97 4.26 1.97 4.26 1.96 2.815 1.96 2.815 1.84 4.38 1.84 4.38 1.85 4.675 1.85 4.675 0.8 4.465 0.8 4.465 0.68 4.795 0.68 ;
      POLYGON 4.315 1.34 3.555 1.34 3.555 0.94 3.675 0.94 3.675 1.22 4.315 1.22 ;
      POLYGON 3.495 1.72 2.695 1.72 2.695 1.76 0.615 1.76 0.615 1 0.735 1 0.735 1.64 2.575 1.64 2.575 1.6 3.315 1.6 3.315 0.88 3.175 0.88 3.175 0.58 3.055 0.58 3.055 0.46 3.295 0.46 3.295 0.76 3.435 0.76 3.435 1.46 3.495 1.46 ;
      POLYGON 1.075 1.17 0.955 1.17 0.955 0.88 0.495 0.88 0.495 1.46 0.255 1.46 0.255 1.99 0.135 1.99 0.135 1.34 0.375 1.34 0.375 0.59 0.495 0.59 0.495 0.76 1.075 0.76 ;
  END
END DLY4X4

MACRO CLKXOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X8 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.365 0.96 3.485 1.36 ;
        RECT 3.205 0.94 3.465 1.165 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.255 1.11 5.495 1.23 ;
        RECT 5.29 1.11 5.44 1.435 ;
        RECT 4.675 1.04 5.41 1.16 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.725 1.41 2.845 2.21 ;
        RECT 2.595 0.715 2.835 0.835 ;
        RECT 2.545 1.41 2.845 1.53 ;
        RECT 0.135 0.76 2.715 0.88 ;
        RECT 0.36 1.29 2.665 1.41 ;
        RECT 1.885 1.29 2.005 2.21 ;
        RECT 1.755 0.71 1.995 0.88 ;
        RECT 1.045 1.29 1.165 2.21 ;
        RECT 0.915 0.71 1.155 0.88 ;
        RECT 0.36 0.76 0.51 1.145 ;
        RECT 0.205 1.41 0.48 1.53 ;
        RECT 0.36 0.76 0.48 1.53 ;
        RECT 0.205 1.41 0.325 2.21 ;
        RECT 0.135 0.64 0.255 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.235 -0.18 5.355 0.68 ;
        RECT 3.015 0.46 3.255 0.58 ;
        RECT 3.015 -0.18 3.135 0.58 ;
        RECT 2.235 -0.18 2.355 0.64 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 4.975 1.76 5.095 2.79 ;
        RECT 3.085 2 3.325 2.15 ;
        RECT 3.085 2 3.205 2.79 ;
        RECT 2.305 1.53 2.425 2.79 ;
        RECT 1.465 1.53 1.585 2.79 ;
        RECT 0.625 1.53 0.745 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.775 0.92 5.735 0.92 5.735 1.675 5.575 1.675 5.575 1.93 5.455 1.93 5.455 1.555 5.615 1.555 5.615 0.92 4.455 0.92 4.455 1.28 4.575 1.28 4.575 1.4 4.335 1.4 4.335 1.04 3.975 1.04 3.975 1.12 3.855 1.12 3.855 0.88 3.975 0.88 3.975 0.92 4.335 0.92 4.335 0.8 5.615 0.8 5.615 0.56 5.655 0.56 5.655 0.44 5.775 0.44 ;
      POLYGON 5.075 1.64 4.035 1.64 4.035 2.01 3.915 2.01 3.915 1.64 3.615 1.64 3.615 0.6 3.875 0.6 3.875 0.72 3.735 0.72 3.735 1.52 4.955 1.52 4.955 1.37 5.075 1.37 ;
      POLYGON 4.455 2.21 4.36 2.21 4.36 2.25 3.445 2.25 3.445 1.88 3.18 1.88 3.18 1.76 2.965 1.76 2.965 1.17 1.935 1.17 1.935 1.05 2.965 1.05 2.965 0.7 3.375 0.7 3.375 0.36 4.235 0.36 4.235 0.68 4.115 0.68 4.115 0.48 3.495 0.48 3.495 0.82 3.085 0.82 3.085 1.64 3.3 1.64 3.3 1.76 3.565 1.76 3.565 2.13 4.24 2.13 4.24 2.09 4.335 2.09 4.335 1.76 4.455 1.76 ;
  END
END CLKXOR2X8

MACRO OR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X8 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.055 1.635 1.175 ;
        RECT 0.36 1.175 0.56 1.295 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.295 1.015 1.415 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.295 0.8 1.725 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.695 0.715 4.935 0.835 ;
        RECT 2.295 0.765 4.815 0.885 ;
        RECT 4.615 1.47 4.735 2.21 ;
        RECT 4.435 1.47 4.735 1.59 ;
        RECT 4.435 1.275 4.555 1.59 ;
        RECT 2.095 1.275 4.555 1.395 ;
        RECT 3.935 0.765 4.28 1.145 ;
        RECT 3.935 0.765 4.055 1.395 ;
        RECT 3.915 0.645 4.035 0.885 ;
        RECT 3.775 1.275 3.895 2.21 ;
        RECT 3.015 0.715 3.255 0.885 ;
        RECT 2.935 1.275 3.055 2.21 ;
        RECT 2.175 0.715 2.415 0.835 ;
        RECT 2.095 1.275 2.215 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 4.335 -0.18 4.455 0.645 ;
        RECT 3.495 -0.18 3.615 0.645 ;
        RECT 2.655 -0.18 2.775 0.645 ;
        RECT 1.815 -0.18 1.935 0.695 ;
        RECT 0.975 -0.18 1.095 0.695 ;
        RECT 0.135 -0.18 0.255 0.695 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.195 1.515 4.315 2.79 ;
        RECT 3.355 1.515 3.475 2.79 ;
        RECT 2.515 1.515 2.635 2.79 ;
        RECT 1.675 1.555 1.795 2.79 ;
        RECT 0.335 1.555 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.815 1.155 1.875 1.155 1.875 1.415 1.255 1.415 1.255 1.675 1.095 1.675 1.095 2.205 0.975 2.205 0.975 1.555 1.135 1.555 1.135 1.295 1.755 1.295 1.755 0.935 0.555 0.935 0.555 0.645 0.675 0.645 0.675 0.815 1.395 0.815 1.395 0.645 1.515 0.645 1.515 0.815 1.875 0.815 1.875 1.035 3.815 1.035 ;
  END
END OR2X8

MACRO DFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFXL 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.03 1.155 2.305 1.38 ;
        RECT 1.925 1.12 2.185 1.315 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.395 1.48 6.695 1.73 ;
        RECT 6.395 1.48 6.655 1.75 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 1.3 0.255 1.58 ;
        RECT 0.135 0.68 0.255 0.94 ;
        RECT 0.115 0.82 0.235 1.42 ;
        RECT 0.07 0.885 0.235 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.38 1.565 1.62 ;
        RECT 1.365 0.68 1.485 0.96 ;
        RECT 1.325 0.84 1.445 1.62 ;
        RECT 1.23 1.465 1.38 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.515 0.67 6.755 0.79 ;
        RECT 6.635 -0.18 6.755 0.79 ;
        RECT 5.015 0.57 5.255 0.69 ;
        RECT 5.135 -0.18 5.255 0.69 ;
        RECT 3.095 -0.18 3.215 0.86 ;
        RECT 1.805 -0.18 1.925 0.4 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.595 1.87 6.715 2.79 ;
        RECT 4.955 2.29 5.195 2.79 ;
        RECT 3.175 2.29 3.415 2.79 ;
        RECT 1.865 1.5 1.985 2.79 ;
        RECT 0.555 1.46 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.175 1.51 7.135 1.51 7.135 1.99 7.015 1.99 7.015 1.39 7.055 1.39 7.055 1.03 6.275 1.03 6.275 0.5 5.595 0.5 5.595 0.93 4.775 0.93 4.775 0.5 4.415 0.5 4.415 1.12 4.295 1.12 4.295 1.33 3.775 1.33 3.775 1.45 3.655 1.45 3.655 1.21 4.175 1.21 4.175 1 4.295 1 4.295 0.38 4.895 0.38 4.895 0.81 5.475 0.81 5.475 0.38 5.575 0.38 5.575 0.36 5.815 0.36 5.815 0.38 6.395 0.38 6.395 0.91 7.055 0.91 7.055 0.62 7.175 0.62 ;
      POLYGON 6.935 1.27 6.815 1.27 6.815 1.36 6.275 1.36 6.275 1.4 6.075 1.4 6.075 2.23 5.315 2.23 5.315 2.17 4.355 2.17 4.355 2.23 3.61 2.23 3.61 2.17 2.285 2.17 2.285 1.5 2.425 1.5 2.425 1 2.285 1 2.285 0.68 2.405 0.68 2.405 0.88 2.545 0.88 2.545 1.62 2.405 1.62 2.405 2.05 3.73 2.05 3.73 2.11 4.235 2.11 4.235 1.61 4.175 1.61 4.175 1.49 4.415 1.49 4.415 1.61 4.355 1.61 4.355 2.05 5.435 2.05 5.435 2.11 5.955 2.11 5.955 1.61 5.515 1.61 5.515 1.49 5.955 1.49 5.955 1.24 6.155 1.24 6.155 1.16 6.275 1.16 6.275 1.24 6.695 1.24 6.695 1.15 6.935 1.15 ;
      POLYGON 5.995 0.86 5.835 0.86 5.835 1.37 5.395 1.37 5.395 1.73 5.835 1.73 5.835 1.99 5.715 1.99 5.715 1.85 5.275 1.85 5.275 1.53 4.915 1.53 4.915 1.65 4.795 1.65 4.795 1.41 5.275 1.41 5.275 1.25 5.715 1.25 5.715 0.74 5.875 0.74 5.875 0.62 5.995 0.62 ;
      POLYGON 5.155 1.29 4.655 1.29 4.655 1.81 4.715 1.81 4.715 1.93 4.475 1.93 4.475 1.81 4.535 1.81 4.535 0.62 4.655 0.62 4.655 1.17 5.035 1.17 5.035 1.05 5.155 1.05 ;
      POLYGON 4.175 0.8 3.79 0.8 3.79 1.09 3.535 1.09 3.535 1.57 4.055 1.57 4.055 1.99 3.935 1.99 3.935 1.69 3.415 1.69 3.415 1.65 3.015 1.65 3.015 1.41 3.135 1.41 3.135 1.53 3.415 1.53 3.415 0.97 3.67 0.97 3.67 0.68 4.175 0.68 ;
      POLYGON 3.295 1.22 2.895 1.22 2.895 1.81 2.935 1.81 2.935 1.93 2.695 1.93 2.695 1.81 2.775 1.81 2.775 0.86 2.675 0.86 2.675 0.56 2.165 0.56 2.165 1 1.805 1 1.805 1.2 1.565 1.2 1.565 1.08 1.685 1.08 1.685 0.88 2.045 0.88 2.045 0.44 2.795 0.44 2.795 0.74 2.895 0.74 2.895 1.1 3.175 1.1 3.175 0.98 3.295 0.98 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.18 0.355 1.18 0.355 1.06 0.975 1.06 0.975 0.68 1.095 0.68 ;
  END
END DFFXL

MACRO OAI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X4 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.465 ;
        RECT 0.375 1.01 0.495 1.495 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.02 0.835 1.4 ;
        RECT 0.65 1.065 0.8 1.435 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.025 1.28 8.265 1.4 ;
        RECT 8.025 1.28 8.145 1.59 ;
        RECT 5.575 1.47 8.145 1.59 ;
        RECT 6.555 1.3 6.795 1.59 ;
        RECT 5.525 1.52 5.785 1.67 ;
        RECT 5.575 1.28 5.695 1.67 ;
        RECT 5.425 1.28 5.695 1.4 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.174 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.4028 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 0.94 6.075 1.17 ;
        RECT 5.845 0.94 5.965 1.35 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.965 0.46 8.205 0.58 ;
        RECT 6.375 0.41 8.085 0.53 ;
        RECT 5.985 1.71 7.785 1.83 ;
        RECT 7.125 0.41 7.365 0.58 ;
        RECT 6.225 0.46 6.525 0.58 ;
        RECT 5.185 0.7 6.345 0.82 ;
        RECT 6.225 0.46 6.345 0.82 ;
        RECT 5.985 1.71 6.105 2.01 ;
        RECT 5.185 1.79 6.105 1.91 ;
        RECT 5.445 0.65 5.685 0.82 ;
        RECT 2.645 1.69 5.305 1.81 ;
        RECT 5.185 0.7 5.305 1.91 ;
        RECT 4.945 1.52 5.305 1.81 ;
        RECT 4.125 1.56 4.245 2.01 ;
        RECT 2.645 1.69 2.765 2.01 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 4.545 -0.18 4.785 0.34 ;
        RECT 3.645 0.46 3.885 0.58 ;
        RECT 3.645 -0.18 3.765 0.58 ;
        RECT 2.805 0.46 3.045 0.58 ;
        RECT 2.805 -0.18 2.925 0.58 ;
        RECT 2.025 -0.18 2.145 0.64 ;
        RECT 0.555 -0.18 0.675 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 8.245 2.19 8.485 2.31 ;
        RECT 8.245 2.19 8.365 2.79 ;
        RECT 6.755 2.19 6.995 2.31 ;
        RECT 6.755 2.19 6.875 2.79 ;
        RECT 5.085 2.27 5.325 2.79 ;
        RECT 3.285 2.17 3.525 2.29 ;
        RECT 3.285 2.17 3.405 2.79 ;
        RECT 2.005 1.93 2.125 2.79 ;
        RECT 0.555 1.615 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.565 0.83 8.505 0.83 8.505 2.07 6.635 2.07 6.635 2.25 5.72 2.25 5.72 2.15 4.78 2.15 4.78 2.25 3.645 2.25 3.645 2.05 3.16 2.05 3.16 2.25 2.245 2.25 2.245 1.81 1.305 1.81 1.305 1.08 1.425 1.08 1.425 0.65 1.665 0.65 1.665 0.77 1.545 0.77 1.545 1.08 2.025 1.08 2.025 1.21 2.505 1.21 2.505 0.83 2.445 0.83 2.445 0.59 2.565 0.59 2.565 0.7 3.285 0.7 3.285 0.59 3.405 0.59 3.405 0.7 4.125 0.7 4.125 0.59 4.245 0.59 4.245 0.7 4.88 0.7 4.88 0.46 5.205 0.46 5.205 0.41 5.985 0.41 5.985 0.46 6.105 0.46 6.105 0.58 5.865 0.58 5.865 0.53 5.325 0.53 5.325 0.58 5 0.58 5 0.82 4.245 0.82 4.245 0.83 4.125 0.83 4.125 0.82 3.405 0.82 3.405 0.83 3.285 0.83 3.285 0.82 2.625 0.82 2.625 1.33 1.905 1.33 1.905 1.2 1.425 1.2 1.425 1.69 2.365 1.69 2.365 2.13 3.04 2.13 3.04 1.93 3.765 1.93 3.765 2.13 4.66 2.13 4.66 2.03 5.84 2.03 5.84 2.13 6.515 2.13 6.515 1.95 8.385 1.95 8.385 0.83 6.825 0.83 6.825 0.77 6.705 0.77 6.705 0.65 6.945 0.65 6.945 0.71 7.545 0.71 7.545 0.65 7.785 0.65 7.785 0.71 8.445 0.71 8.445 0.59 8.565 0.59 ;
      POLYGON 7.535 1.18 6.435 1.18 6.435 1.29 6.195 1.29 6.195 1.17 6.315 1.17 6.315 1.06 7.535 1.06 ;
      POLYGON 5.005 1.4 3.325 1.4 3.325 1.57 1.665 1.57 1.665 1.44 1.545 1.44 1.545 1.32 1.785 1.32 1.785 1.45 3.085 1.45 3.085 1.28 5.005 1.28 ;
      RECT 2.745 1 4.025 1.12 ;
      POLYGON 2.385 1.09 2.145 1.09 2.145 0.96 1.785 0.96 1.785 0.48 0.915 0.48 0.915 0.89 0.24 0.89 0.24 1.585 0.255 1.585 0.255 2.21 0.135 2.21 0.135 1.705 0.12 1.705 0.12 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.77 0.795 0.77 0.795 0.36 1.905 0.36 1.905 0.84 2.265 0.84 2.265 0.97 2.385 0.97 ;
      POLYGON 1.185 1.25 1.155 1.25 1.155 1.68 1.095 1.68 1.095 2.21 0.975 2.21 0.975 1.56 1.035 1.56 1.035 0.6 1.155 0.6 1.155 1.01 1.185 1.01 ;
  END
END OAI2BB2X4

MACRO EDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX1 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.8 1.435 ;
        RECT 0.435 1.175 0.8 1.355 ;
        RECT 0.435 1.115 0.555 1.355 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.105 1.13 6.385 1.37 ;
        RECT 6.105 1.13 6.365 1.39 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.545 1.175 6.89 1.435 ;
        RECT 5.565 1.51 6.665 1.63 ;
        RECT 6.545 1.175 6.665 1.63 ;
        RECT 5.185 2.13 5.745 2.25 ;
        RECT 5.625 1.51 5.745 2.25 ;
        RECT 5.565 0.92 5.685 1.63 ;
        RECT 5.445 0.92 5.685 1.04 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.35 0.885 7.47 1.99 ;
        RECT 7.315 0.68 7.435 1.025 ;
        RECT 7.32 0.885 7.47 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.025 0.59 9.145 2.21 ;
        RECT 8.77 1.175 9.145 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 8.545 -0.18 8.665 0.53 ;
        RECT 7.83 -0.18 7.95 0.4 ;
        RECT 6.025 0.41 6.265 0.53 ;
        RECT 6.025 -0.18 6.145 0.53 ;
        RECT 4.485 -0.18 4.605 0.77 ;
        RECT 2.585 0.35 2.825 0.47 ;
        RECT 2.705 -0.18 2.825 0.47 ;
        RECT 0.595 -0.18 0.715 0.695 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 8.605 1.73 8.725 2.79 ;
        RECT 7.77 1.36 7.89 2.79 ;
        RECT 6.365 1.75 6.485 2.79 ;
        RECT 4.365 2.13 4.605 2.25 ;
        RECT 4.365 2.13 4.485 2.79 ;
        RECT 2.585 1.91 2.825 2.03 ;
        RECT 2.585 1.91 2.705 2.79 ;
        RECT 0.595 1.555 0.715 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.65 1.18 8.395 1.18 8.395 1.3 8.37 1.3 8.37 1.58 8.25 1.58 8.25 1.18 8.275 1.18 8.275 0.68 8.395 0.68 8.395 1.06 8.65 1.06 ;
      POLYGON 7.71 1.24 7.59 1.24 7.59 0.48 6.505 0.48 6.505 0.77 5.785 0.77 5.785 0.48 5.025 0.48 5.025 0.77 5.045 0.77 5.045 1.51 4.965 1.51 4.965 1.65 5.085 1.65 5.085 1.77 4.845 1.77 4.845 1.51 4.365 1.51 4.365 1.27 4.485 1.27 4.485 1.39 4.925 1.39 4.925 0.89 4.905 0.89 4.905 0.36 5.905 0.36 5.905 0.65 6.385 0.65 6.385 0.36 7.71 0.36 ;
      POLYGON 7.13 1.675 6.905 1.675 6.905 1.87 6.785 1.87 6.785 1.555 7.01 1.555 7.01 1.01 5.985 1.01 5.985 1.39 5.865 1.39 5.865 0.89 7.01 0.89 7.01 0.72 6.625 0.72 6.625 0.6 7.13 0.6 ;
      POLYGON 5.565 0.72 5.325 0.72 5.325 1.75 5.505 1.75 5.505 2.01 4.18 2.01 4.18 2.11 2.945 2.11 2.945 1.79 2.465 1.79 2.465 2.11 1.525 2.11 1.525 1.87 1.345 1.87 1.345 0.74 1.405 0.74 1.405 0.62 1.525 0.62 1.525 0.86 1.465 0.86 1.465 1.75 1.645 1.75 1.645 1.99 2.345 1.99 2.345 1.67 3.065 1.67 3.065 1.99 4.06 1.99 4.06 1.89 5.205 1.89 5.205 0.6 5.565 0.6 ;
      POLYGON 4.805 1.13 4.245 1.13 4.245 1.77 3.905 1.77 3.905 1.81 3.665 1.81 3.665 1.69 3.785 1.69 3.785 1.65 4.125 1.65 4.125 1.13 3.665 1.13 3.665 0.62 3.785 0.62 3.785 1.01 4.805 1.01 ;
      POLYGON 4.005 1.53 3.885 1.53 3.885 1.41 3.425 1.41 3.425 1.31 3.345 1.31 3.345 1.07 3.425 1.07 3.425 0.5 3.065 0.5 3.065 0.71 2.345 0.71 2.345 0.5 1.765 0.5 1.765 1.37 1.825 1.37 1.825 1.49 1.585 1.49 1.585 1.37 1.645 1.37 1.645 0.5 1.135 0.5 1.135 1.675 1.015 1.675 1.015 0.38 2.025 0.38 2.025 0.36 2.265 0.36 2.265 0.38 2.465 0.38 2.465 0.59 2.945 0.59 2.945 0.38 3.545 0.38 3.545 1.29 4.005 1.29 ;
      POLYGON 3.305 0.95 3.225 0.95 3.225 1.43 3.305 1.43 3.305 1.87 3.185 1.87 3.185 1.55 2.505 1.55 2.505 1.49 2.385 1.49 2.385 1.37 2.625 1.37 2.625 1.43 3.105 1.43 3.105 0.83 3.185 0.83 3.185 0.62 3.305 0.62 ;
      POLYGON 2.985 1.22 2.125 1.22 2.125 1.75 2.065 1.75 2.065 1.87 1.945 1.87 1.945 1.63 2.005 1.63 2.005 0.8 1.885 0.8 1.885 0.68 2.125 0.68 2.125 1.1 2.985 1.1 ;
      POLYGON 0.895 1.055 0.775 1.055 0.775 0.995 0.295 0.995 0.295 1.675 0.175 1.675 0.175 0.455 0.295 0.455 0.295 0.875 0.775 0.875 0.775 0.815 0.895 0.815 ;
  END
END EDFFX1

MACRO HOLDX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HOLDX1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.485 0.68 1.605 1.6 ;
        RECT 0.405 1.36 1.605 1.48 ;
        RECT 1.23 1.175 1.605 1.48 ;
        RECT 0.405 1.02 0.525 1.48 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.885 1.24 0.765 1.24 0.765 0.9 0.255 0.9 0.255 1.99 0.135 1.99 0.135 0.66 0.255 0.66 0.255 0.78 0.885 0.78 ;
  END
END HOLDX1

MACRO OAI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X4 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.73 1.23 8.43 1.35 ;
        RECT 7.845 1.23 8.105 1.38 ;
    END
  END C0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.105 1.23 6.365 1.38 ;
        RECT 6.105 1.06 6.33 1.38 ;
        RECT 4.99 1.06 6.33 1.18 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 1.01 2.94 1.13 ;
        RECT 1.175 1.23 1.435 1.38 ;
        RECT 1.195 1.01 1.435 1.38 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.74 1.175 6.89 1.435 ;
        RECT 4.31 1.5 6.86 1.62 ;
        RECT 6.74 1.175 6.86 1.62 ;
        RECT 5.68 1.3 5.92 1.62 ;
        RECT 4.31 1.22 4.43 1.62 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.5 3.54 1.62 ;
        RECT 3.42 1.24 3.54 1.62 ;
        RECT 2.02 1.25 2.14 1.62 ;
        RECT 0.68 1.175 0.8 1.62 ;
        RECT 0.65 1.175 0.8 1.435 ;
        RECT 0.56 1.3 0.8 1.42 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.55 0.885 8.92 1.145 ;
        RECT 7.73 0.77 8.69 0.89 ;
        RECT 8.57 0.6 8.69 1.145 ;
        RECT 1.12 1.74 8.67 1.86 ;
        RECT 8.37 1.56 8.67 1.86 ;
        RECT 8.55 0.72 8.67 1.86 ;
        RECT 8.37 1.56 8.49 2.21 ;
        RECT 7.73 0.6 7.85 0.89 ;
        RECT 7.53 1.56 7.65 2.21 ;
        RECT 6.24 1.74 6.36 2.21 ;
        RECT 4.96 1.74 5.08 2.21 ;
        RECT 2.92 1.74 3.04 2.21 ;
        RECT 1.12 1.74 1.24 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 3.56 -0.18 3.68 0.65 ;
        RECT 2.72 -0.18 2.84 0.65 ;
        RECT 1.88 -0.18 2 0.65 ;
        RECT 1.04 -0.18 1.16 0.65 ;
        RECT 0.2 -0.18 0.32 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 8.79 1.56 8.91 2.79 ;
        RECT 7.89 1.98 8.13 2.15 ;
        RECT 7.89 1.98 8.01 2.79 ;
        RECT 7.05 1.98 7.29 2.15 ;
        RECT 7.05 1.98 7.17 2.79 ;
        RECT 5.54 1.98 5.78 2.15 ;
        RECT 5.54 1.98 5.66 2.79 ;
        RECT 3.5 1.98 3.74 2.15 ;
        RECT 3.5 1.98 3.62 2.79 ;
        RECT 1.7 1.98 1.94 2.15 ;
        RECT 1.7 1.98 1.82 2.79 ;
        RECT 0.48 1.74 0.6 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.11 0.65 8.99 0.65 8.99 0.48 8.27 0.48 8.27 0.65 8.15 0.65 8.15 0.48 7.43 0.48 7.43 0.65 7.31 0.65 7.31 0.48 6.59 0.48 6.59 0.65 6.47 0.65 6.47 0.48 5.75 0.48 5.75 0.65 5.63 0.65 5.63 0.48 4.91 0.48 4.91 0.65 4.79 0.65 4.79 0.48 4.07 0.48 4.07 0.65 3.95 0.65 3.95 0.36 9.11 0.36 ;
      POLYGON 7.07 0.78 6.95 0.78 6.95 0.89 0.62 0.89 0.62 0.6 0.74 0.6 0.74 0.77 1.46 0.77 1.46 0.6 1.58 0.6 1.58 0.77 2.3 0.77 2.3 0.6 2.42 0.6 2.42 0.77 3.14 0.77 3.14 0.6 3.26 0.6 3.26 0.77 4.37 0.77 4.37 0.6 4.49 0.6 4.49 0.77 5.21 0.77 5.21 0.6 5.33 0.6 5.33 0.77 6.05 0.77 6.05 0.6 6.17 0.6 6.17 0.77 6.83 0.77 6.83 0.66 7.07 0.66 ;
  END
END OAI221X4

MACRO ANTENNA
  CLASS CORE ANTENNACELL ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.116 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.185 0.3 0.685 2.31 ;
    END
  END A
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
    END
  END VDD
END ANTENNA

MACRO OAI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X1 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 1.18 0.565 1.67 ;
        RECT 0.305 1.18 0.565 1.4 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.52 1.145 1.705 ;
        RECT 0.885 1.33 1.005 1.705 ;
    END
  END A0N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.15 3.12 1.435 ;
        RECT 2.855 1.1 2.975 1.37 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 0.885 3.7 1.2 ;
        RECT 3.48 1.08 3.6 1.39 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.475 1.555 3.36 1.675 ;
        RECT 3.24 0.8 3.36 1.675 ;
        RECT 3.095 0.8 3.36 0.92 ;
        RECT 3.095 0.68 3.215 0.92 ;
        RECT 2.675 1.53 2.795 2.18 ;
        RECT 2.335 1.53 2.795 1.67 ;
        RECT 2.335 1.52 2.595 1.67 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 2.195 0.55 2.435 0.67 ;
        RECT 2.195 -0.18 2.315 0.67 ;
        RECT 0.685 -0.18 0.805 0.82 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.48 1.53 3.6 2.79 ;
        RECT 2.035 1.53 2.155 2.79 ;
        RECT 0.625 1.825 0.745 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.635 0.73 3.515 0.73 3.515 0.61 3.385 0.61 3.385 0.56 2.975 0.56 2.975 0.91 1.835 0.91 1.835 0.67 1.955 0.67 1.955 0.79 2.615 0.79 2.615 0.74 2.855 0.74 2.855 0.44 3.505 0.44 3.505 0.49 3.635 0.49 ;
      POLYGON 2.695 1.2 2.455 1.2 2.455 1.15 1.595 1.15 1.595 0.48 1.045 0.48 1.045 1.06 0.185 1.06 0.185 1.705 0.325 1.705 0.325 1.945 0.205 1.945 0.205 1.825 0.065 1.825 0.065 0.72 0.205 0.72 0.205 0.6 0.325 0.6 0.325 0.94 0.925 0.94 0.925 0.36 1.715 0.36 1.715 1.03 2.575 1.03 2.575 1.08 2.695 1.08 ;
      POLYGON 2.155 1.39 1.385 1.39 1.385 1.945 1.165 1.945 1.165 2.065 1.045 2.065 1.045 1.825 1.265 1.825 1.265 0.84 1.165 0.84 1.165 0.6 1.285 0.6 1.285 0.72 1.385 0.72 1.385 1.27 2.155 1.27 ;
  END
END OAI2BB2X1

MACRO CLKINVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX1 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.795 0.24 1.22 ;
        RECT 0.07 0.795 0.24 1.2 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.625 0.675 1.99 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
        RECT 0.135 -0.18 0.255 0.675 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
END CLKINVX1

MACRO SDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX2 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.465 1.335 1.585 ;
        RECT 1.215 1.345 1.335 1.585 ;
        RECT 0.94 1.465 1.09 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.485 0.96 6.68 1.2 ;
        RECT 6.45 0.885 6.675 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.9 1.025 8.06 1.48 ;
        RECT 7.94 1 8.06 1.48 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 1.23 8.685 1.38 ;
        RECT 8.425 1.07 8.545 1.38 ;
        RECT 8.34 0.76 8.46 1.19 ;
        RECT 8.22 1.07 8.545 1.19 ;
        RECT 7.3 0.76 8.46 0.88 ;
        RECT 7.54 0.76 7.78 1.09 ;
        RECT 7.04 1 7.42 1.12 ;
        RECT 7.3 0.76 7.42 1.12 ;
        RECT 7.04 1 7.16 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.68 0.675 2.205 ;
        RECT 0.36 1.175 0.675 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.1 -0.18 8.22 0.64 ;
        RECT 6.82 -0.18 6.94 0.64 ;
        RECT 4.43 0.38 4.67 0.5 ;
        RECT 4.55 -0.18 4.67 0.5 ;
        RECT 2.57 -0.18 2.69 0.68 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 7.94 1.84 8.06 2.79 ;
        RECT 6.56 1.56 6.68 2.79 ;
        RECT 4.43 2.06 4.67 2.18 ;
        RECT 4.43 2.06 4.55 2.79 ;
        RECT 2.31 2.06 2.43 2.79 ;
        RECT 0.975 1.845 1.095 2.79 ;
        RECT 0.135 1.555 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.925 1.72 8.54 1.72 8.54 1.84 8.42 1.84 8.42 1.72 7.44 1.72 7.44 1.24 7.56 1.24 7.56 1.6 8.805 1.6 8.805 0.95 8.58 0.95 8.58 0.59 8.7 0.59 8.7 0.83 8.925 0.83 ;
      POLYGON 7.58 0.64 7.18 0.64 7.18 0.88 6.92 0.88 6.92 1.56 7.32 1.56 7.32 2.21 7.2 2.21 7.2 1.68 6.8 1.68 6.8 1.44 5.99 1.44 5.99 1.58 5.95 1.58 5.95 1.7 5.83 1.7 5.83 1.46 5.87 1.46 5.87 0.72 5.83 0.72 5.83 0.6 6.07 0.6 6.07 0.72 5.99 0.72 5.99 1.32 6.8 1.32 6.8 0.76 7.06 0.76 7.06 0.52 7.46 0.52 7.46 0.4 7.58 0.4 ;
      POLYGON 6.46 0.66 6.34 0.66 6.34 0.48 5.71 0.48 5.71 1.1 5.75 1.1 5.75 1.34 5.71 1.34 5.71 1.91 6.26 1.91 6.26 2.03 5.59 2.03 5.59 0.48 5.11 0.48 5.11 0.92 5.23 0.92 5.23 1.04 4.99 1.04 4.99 0.74 4.19 0.74 4.19 0.48 3.71 0.48 3.71 0.98 3.57 0.98 3.57 1.26 2.99 1.26 2.99 1.38 2.87 1.38 2.87 1.14 3.45 1.14 3.45 0.86 3.59 0.86 3.59 0.36 4.31 0.36 4.31 0.62 4.99 0.62 4.99 0.36 6.46 0.36 ;
      POLYGON 5.47 1.98 5.35 1.98 5.35 1.3 4.29 1.3 4.29 1.18 5.35 1.18 5.35 0.72 5.23 0.72 5.23 0.6 5.47 0.6 ;
      POLYGON 5.25 2.24 5.01 2.24 5.01 1.94 3.89 1.94 3.89 2.22 2.71 2.22 2.71 1.94 2.035 1.94 2.035 1.965 1.515 1.965 1.515 2.085 1.395 2.085 1.395 1.845 1.455 1.845 1.455 0.68 1.575 0.68 1.575 1.845 1.915 1.845 1.915 1.82 2.83 1.82 2.83 2.1 3.77 2.1 3.77 1.22 3.81 1.22 3.81 1.1 3.93 1.1 3.93 1.34 3.89 1.34 3.89 1.82 5.13 1.82 5.13 2.12 5.25 2.12 ;
      POLYGON 4.87 1.06 4.17 1.06 4.17 1.58 4.13 1.58 4.13 1.7 4.01 1.7 4.01 1.46 4.05 1.46 4.05 0.98 3.83 0.98 3.83 0.6 4.07 0.6 4.07 0.86 4.17 0.86 4.17 0.94 4.87 0.94 ;
      POLYGON 3.47 0.72 2.93 0.72 2.93 1.02 2.75 1.02 2.75 1.5 3.11 1.5 3.11 1.46 3.23 1.46 3.23 1.98 3.11 1.98 3.11 1.62 2.07 1.62 2.07 1.34 2.05 1.34 2.05 1.1 2.19 1.1 2.19 1.5 2.63 1.5 2.63 0.9 2.81 0.9 2.81 0.6 3.47 0.6 ;
      POLYGON 2.51 1.38 2.39 1.38 2.39 0.98 1.93 0.98 1.93 1.46 1.95 1.46 1.95 1.7 1.83 1.7 1.83 1.58 1.81 1.58 1.81 0.56 1.335 0.56 1.335 1.18 0.795 1.18 0.795 1.06 1.215 1.06 1.215 0.44 2.27 0.44 2.27 0.86 2.51 0.86 ;
  END
END SDFFHQX2

MACRO SDFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX8 0 0 ;
  SIZE 16.24 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.32 2.775 2.185 ;
        RECT 2.655 0.68 2.775 0.96 ;
        RECT 0.07 1.2 2.755 1.32 ;
        RECT 2.635 0.84 2.755 1.44 ;
        RECT 1.815 0.68 1.935 2.185 ;
        RECT 0.975 0.68 1.095 2.18 ;
        RECT 0.135 0.68 0.255 2.18 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 1.17 5.245 1.39 ;
        RECT 4.945 1.17 5.205 1.41 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.095 2.13 10.315 2.25 ;
        RECT 9.095 1.7 9.215 2.25 ;
        RECT 8.495 1.7 9.215 1.82 ;
        RECT 7.535 2.13 8.615 2.25 ;
        RECT 8.495 1.7 8.615 2.25 ;
        RECT 7.295 2.08 7.655 2.2 ;
        RECT 7.295 1.42 7.415 2.2 ;
        RECT 5.61 1.42 7.415 1.54 ;
        RECT 5.58 1.21 5.805 1.435 ;
        RECT 5.58 1.175 5.73 1.435 ;
        RECT 5.565 1.21 5.805 1.33 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.415 0.96 13.535 1.2 ;
        RECT 13.065 0.96 13.535 1.09 ;
        RECT 13.065 0.94 13.325 1.09 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.755 0.755 13.875 1.18 ;
        RECT 13.7 1.035 13.85 1.44 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.935 1.22 15.355 1.44 ;
        RECT 15.095 1.2 15.355 1.44 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.73 1.175 15.88 1.435 ;
        RECT 15.555 0.96 15.85 1.2 ;
        RECT 14.235 0.96 15.85 1.08 ;
        RECT 14.735 0.96 14.975 1.1 ;
        RECT 14.235 0.96 14.355 1.44 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 16.24 0.18 ;
        RECT 15.295 -0.18 15.415 0.84 ;
        RECT 13.775 -0.18 14.015 0.32 ;
        RECT 12.725 -0.18 12.965 0.32 ;
        RECT 10.615 -0.18 10.735 0.68 ;
        RECT 5.265 0.69 5.505 0.81 ;
        RECT 5.385 -0.18 5.505 0.81 ;
        RECT 3.915 -0.18 4.035 0.665 ;
        RECT 3.075 -0.18 3.195 0.665 ;
        RECT 2.235 -0.18 2.355 0.67 ;
        RECT 1.395 -0.18 1.515 0.67 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 16.24 2.79 ;
        RECT 15.075 1.8 15.195 2.79 ;
        RECT 13.755 1.56 13.875 2.79 ;
        RECT 12.845 1.56 12.965 2.79 ;
        RECT 10.475 1.88 10.715 2 ;
        RECT 10.475 1.88 10.595 2.79 ;
        RECT 8.855 1.94 8.975 2.79 ;
        RECT 8.735 1.94 8.975 2.06 ;
        RECT 6.605 1.9 6.845 2.02 ;
        RECT 6.605 1.9 6.725 2.79 ;
        RECT 5.205 1.9 5.445 2.02 ;
        RECT 5.205 1.9 5.325 2.79 ;
        RECT 3.915 1.535 4.035 2.79 ;
        RECT 3.075 1.535 3.195 2.79 ;
        RECT 2.235 1.44 2.355 2.79 ;
        RECT 1.395 1.44 1.515 2.79 ;
        RECT 0.555 1.44 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 16.12 1.98 15.435 1.98 15.435 1.86 16 1.86 16 1.68 14.635 1.68 14.635 1.42 14.515 1.42 14.515 1.3 14.755 1.3 14.755 1.56 16 1.56 16 0.84 15.715 0.84 15.715 0.6 15.835 0.6 15.835 0.72 16.12 0.72 ;
      POLYGON 14.715 0.635 14.115 0.635 14.115 1.56 14.515 1.56 14.515 2.21 14.395 2.21 14.395 1.68 13.995 1.68 13.995 0.635 13.73 0.635 13.73 0.56 11.795 0.56 11.795 1 12.135 1 12.135 1.58 12.155 1.58 12.155 1.77 11.915 1.77 11.915 1.58 12.015 1.58 12.015 1.12 11.675 1.12 11.675 0.44 13.85 0.44 13.85 0.515 14.715 0.515 ;
      POLYGON 13.515 1.74 13.275 1.74 13.275 1.44 12.725 1.44 12.725 2.25 10.835 2.25 10.835 1.76 10.355 1.76 10.355 2.01 9.335 2.01 9.335 1.58 8.375 1.58 8.375 2.01 7.775 2.01 7.775 0.98 7.875 0.98 7.875 0.48 7.395 0.48 7.395 1.06 7.155 1.06 7.155 0.94 7.275 0.94 7.275 0.36 7.995 0.36 7.995 1.1 7.895 1.1 7.895 1.89 8.255 1.89 8.255 1.46 9.455 1.46 9.455 1.89 10.235 1.89 10.235 1.64 10.955 1.64 10.955 2.13 12.605 2.13 12.605 0.7 13.195 0.7 13.195 0.68 13.435 0.68 13.435 0.8 13.315 0.8 13.315 0.82 12.725 0.82 12.725 1.32 13.395 1.32 13.395 1.62 13.515 1.62 ;
      POLYGON 12.485 2.01 11.075 2.01 11.075 1.28 11.055 1.28 11.055 1.16 10.575 1.16 10.575 1.28 9.815 1.28 9.815 1.1 8.475 1.1 8.475 1.04 8.355 1.04 8.355 0.92 8.595 0.92 8.595 0.98 9.935 0.98 9.935 1.16 10.455 1.16 10.455 1.04 11.295 1.04 11.295 1.16 11.195 1.16 11.195 1.89 11.675 1.89 11.675 1.36 11.655 1.36 11.655 1.24 11.895 1.24 11.895 1.36 11.795 1.36 11.795 1.89 12.365 1.89 12.365 0.8 12.245 0.8 12.245 0.68 12.485 0.68 ;
      POLYGON 11.555 1.77 11.315 1.77 11.315 1.6 11.415 1.6 11.415 0.78 11.11 0.78 11.11 0.92 10.295 0.92 10.295 1.04 10.055 1.04 10.055 0.92 10.175 0.92 10.175 0.8 10.99 0.8 10.99 0.66 11.255 0.66 11.255 0.54 11.375 0.54 11.375 0.66 11.535 0.66 11.535 1.6 11.555 1.6 ;
      POLYGON 10.935 1.4 10.815 1.4 10.815 1.52 10.115 1.52 10.115 1.77 9.995 1.77 9.995 1.52 9.575 1.52 9.575 1.34 8.135 1.34 8.135 1.77 8.015 1.77 8.015 1.22 8.115 1.22 8.115 0.54 8.235 0.54 8.235 0.68 9.04 0.68 9.04 0.74 9.715 0.74 9.715 0.6 9.955 0.6 9.955 0.72 9.835 0.72 9.835 0.86 8.92 0.86 8.92 0.8 8.235 0.8 8.235 1.22 9.695 1.22 9.695 1.4 10.695 1.4 10.695 1.28 10.935 1.28 ;
      POLYGON 10.315 0.68 10.195 0.68 10.195 0.48 9.535 0.48 9.535 0.62 9.295 0.62 9.295 0.5 9.415 0.5 9.415 0.36 10.315 0.36 ;
      POLYGON 7.755 0.72 7.655 0.72 7.655 1.96 7.535 1.96 7.535 1.3 5.925 1.3 5.925 1.055 5.365 1.055 5.365 1.05 5.025 1.05 5.025 0.495 4.275 0.495 4.275 1.175 4.155 1.175 4.155 0.375 5.145 0.375 5.145 0.93 5.485 0.93 5.485 0.935 6.045 0.935 6.045 1.18 7.535 1.18 7.535 0.72 7.515 0.72 7.515 0.6 7.755 0.6 ;
      POLYGON 7.175 1.96 7.055 1.96 7.055 1.78 5.925 1.78 5.925 1.99 5.805 1.99 5.805 1.66 7.175 1.66 ;
      POLYGON 7.155 0.72 7.035 0.72 7.035 1.055 6.165 1.055 6.165 0.675 6.285 0.675 6.285 0.935 6.915 0.935 6.915 0.6 7.155 0.6 ;
      POLYGON 6.705 0.815 6.585 0.815 6.585 0.555 5.91 0.555 5.91 0.575 5.865 0.575 5.865 0.815 5.745 0.815 5.745 0.455 5.79 0.455 5.79 0.435 6.705 0.435 ;
      POLYGON 6.485 2.25 5.565 2.25 5.565 1.78 5.3 1.78 5.3 1.77 4.785 1.77 4.785 1.65 4.705 1.65 4.705 0.93 4.785 0.93 4.785 0.63 4.905 0.63 4.905 1.05 4.825 1.05 4.825 1.53 4.905 1.53 4.905 1.65 5.42 1.65 5.42 1.66 5.685 1.66 5.685 2.13 6.485 2.13 ;
      POLYGON 5.085 2.25 4.335 2.25 4.335 1.535 4.395 1.535 4.395 1.415 3.615 1.415 3.615 2.185 3.495 2.185 3.495 1.2 2.875 1.2 2.875 1.08 3.495 1.08 3.495 0.615 3.615 0.615 3.615 1.295 4.395 1.295 4.395 0.615 4.515 0.615 4.515 1.655 4.455 1.655 4.455 2.13 5.085 2.13 ;
  END
END SDFFSRHQX8

MACRO CLKXOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.22 1.335 1.46 ;
        RECT 0.885 1.23 1.335 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.18 3.175 1.3 ;
        RECT 2.335 1.18 2.595 1.38 ;
        RECT 2.255 1.14 2.495 1.3 ;
        RECT 1.695 1.34 1.935 1.46 ;
        RECT 1.815 1.18 1.935 1.46 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.74 0.715 2.21 ;
        RECT 0.405 0.74 0.675 0.86 ;
        RECT 0.555 0.62 0.675 0.86 ;
        RECT 0.405 1.74 0.715 1.86 ;
        RECT 0.405 0.74 0.525 1.86 ;
        RECT 0.36 0.885 0.525 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.735 -0.18 2.855 0.78 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.615 1.74 2.735 2.79 ;
        RECT 1.015 2.22 1.255 2.79 ;
        RECT 0.165 1.56 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.415 1.74 3.155 1.74 3.155 1.86 3.035 1.86 3.035 1.62 2.335 1.62 2.335 2.24 2.055 2.24 2.055 2.12 2.215 2.12 2.215 1.5 3.155 1.5 3.155 1.62 3.295 1.62 3.295 0.78 3.155 0.78 3.155 0.54 3.275 0.54 3.275 0.66 3.415 0.66 ;
      POLYGON 2.855 1.06 2.615 1.06 2.615 1.02 1.575 1.02 1.575 1.58 1.675 1.58 1.675 1.86 1.555 1.86 1.555 1.7 1.455 1.7 1.455 0.6 1.695 0.6 1.695 0.72 1.575 0.72 1.575 0.9 2.735 0.9 2.735 0.94 2.855 0.94 ;
      POLYGON 2.215 0.78 2.095 0.78 2.095 0.48 1.335 0.48 1.335 1.1 0.765 1.1 0.765 1.5 0.955 1.5 0.955 1.58 1.14 1.58 1.14 1.98 1.815 1.98 1.815 1.86 1.975 1.86 1.975 1.74 2.095 1.74 2.095 1.98 1.935 1.98 1.935 2.1 1.02 2.1 1.02 1.7 0.835 1.7 0.835 1.62 0.645 1.62 0.645 0.98 1.215 0.98 1.215 0.36 2.215 0.36 ;
  END
END CLKXOR2X2

MACRO TLATNTSCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX8 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.825 0.565 1.09 ;
        RECT 0.325 0.78 0.565 1.09 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.76 1.09 1.23 ;
        RECT 0.925 0.76 1.045 1.26 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.8 1.385 1.26 ;
        RECT 1.23 0.76 1.38 1.195 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.3 1.225 9.42 2.205 ;
        RECT 9.26 0.645 9.38 1.345 ;
        RECT 6.74 1.225 9.42 1.345 ;
        RECT 7.64 0.765 9.38 0.885 ;
        RECT 8.36 0.715 8.6 0.885 ;
        RECT 8.46 1.225 8.58 2.205 ;
        RECT 7.52 0.715 7.76 0.835 ;
        RECT 7.62 1.225 7.74 2.21 ;
        RECT 6.78 0.775 6.9 2.21 ;
        RECT 6.74 0.655 6.86 0.895 ;
        RECT 6.74 1.175 6.9 1.435 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.84 -0.18 8.96 0.645 ;
        RECT 8 -0.18 8.12 0.645 ;
        RECT 7.16 -0.18 7.28 0.645 ;
        RECT 6.32 -0.18 6.44 0.64 ;
        RECT 5.04 -0.18 5.16 0.74 ;
        RECT 3.35 0.41 3.59 0.53 ;
        RECT 3.47 -0.18 3.59 0.53 ;
        RECT 1.08 -0.18 1.2 0.64 ;
        RECT 0.24 -0.18 0.36 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.88 1.465 9 2.79 ;
        RECT 8.04 1.465 8.16 2.79 ;
        RECT 7.2 1.465 7.32 2.79 ;
        RECT 6.36 1.77 6.48 2.79 ;
        RECT 5.52 1.77 5.64 2.79 ;
        RECT 4.66 1.69 4.78 2.79 ;
        RECT 3.25 2 3.37 2.79 ;
        RECT 3.13 2 3.37 2.12 ;
        RECT 0.96 1.62 1.08 2.79 ;
        RECT 0.84 1.62 1.08 1.74 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.62 1.215 6.4 1.215 6.4 1.65 6.06 1.65 6.06 2.21 5.94 2.21 5.94 1.65 5.22 1.65 5.22 2.21 5.1 2.21 5.1 1.53 6.28 1.53 6.28 1.05 5.76 1.05 5.76 0.81 5.68 0.81 5.68 0.57 5.8 0.57 5.8 0.69 5.88 0.69 5.88 0.93 6.62 0.93 ;
      POLYGON 6.16 1.41 5.04 1.41 5.04 1.25 4.3 1.25 4.3 2.01 4.18 2.01 4.18 1.4 3.13 1.4 3.13 1.28 4.18 1.28 4.18 1.13 4.56 1.13 4.56 0.6 4.68 0.6 4.68 1.13 5.16 1.13 5.16 1.29 6.04 1.29 6.04 1.17 6.16 1.17 ;
      POLYGON 5.64 1.17 5.52 1.17 5.52 1.05 5.44 1.05 5.44 0.98 4.8 0.98 4.8 0.48 4.19 0.48 4.19 0.76 4.07 0.76 4.07 1.01 4.06 1.01 4.06 1.16 3.01 1.16 3.01 1.52 3.85 1.52 3.85 1.88 3.97 1.88 3.97 2 3.73 2 3.73 1.64 2.89 1.64 2.89 1.3 2.85 1.3 2.85 1.04 3.94 1.04 3.94 0.89 3.95 0.89 3.95 0.64 4.07 0.64 4.07 0.36 4.92 0.36 4.92 0.86 5.56 0.86 5.56 0.93 5.64 0.93 ;
      POLYGON 4.54 2.25 3.49 2.25 3.49 1.88 2.67 1.88 2.67 2.06 2.55 2.06 2.55 1.94 2.37 1.94 2.37 0.82 2.25 0.82 2.25 0.7 2.49 0.7 2.49 1.76 3.61 1.76 3.61 2.13 4.42 2.13 4.42 1.37 4.54 1.37 ;
      POLYGON 3.95 0.48 3.83 0.48 3.83 0.77 2.73 0.77 2.73 1.64 2.61 1.64 2.61 0.58 2.345 0.58 2.345 0.52 1.625 0.52 1.625 1.5 1.68 1.5 1.68 1.62 1.44 1.62 1.44 1.5 1.505 1.5 1.505 0.64 1.5 0.64 1.5 0.4 2.11 0.4 2.11 0.38 2.35 0.38 2.35 0.4 2.465 0.4 2.465 0.46 2.73 0.46 2.73 0.65 3.71 0.65 3.71 0.36 3.95 0.36 ;
      POLYGON 2.25 2.06 2.13 2.06 2.13 1.94 1.2 1.94 1.2 1.5 0.38 1.5 0.38 1.68 0.26 1.68 0.26 1.38 0.685 1.38 0.685 0.66 0.66 0.66 0.66 0.4 0.78 0.4 0.78 0.54 0.805 0.54 0.805 1.38 1.32 1.38 1.32 1.82 1.89 1.82 1.89 0.64 2.01 0.64 2.01 1.82 2.25 1.82 ;
  END
END TLATNTSCAX8

MACRO XNOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X1 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4014 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.27 1.56 8.51 2.25 ;
        RECT 8.39 0.36 8.51 2.25 ;
        RECT 8.135 0.65 8.51 0.8 ;
        RECT 8.27 0.36 8.51 0.8 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.099 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.07 0.325 1.47 ;
        RECT 0.07 1.175 0.325 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.267 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.84 1.045 1.025 1.375 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 1.35 6.81 1.47 ;
        RECT 6.08 1.23 6.365 1.47 ;
        RECT 6.08 0.905 6.2 1.47 ;
        RECT 5.7 0.905 6.2 1.025 ;
    END
  END C
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.73 2.29 7.97 2.79 ;
        RECT 7.79 1.69 7.91 2.79 ;
        RECT 1.865 2.27 2.105 2.79 ;
        RECT 0.685 2.29 0.925 2.79 ;
        RECT 0.745 1.97 0.865 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.73 -0.18 7.97 0.32 ;
        RECT 7.79 -0.18 7.91 0.67 ;
        RECT 1.865 -0.18 2.105 0.32 ;
        RECT 0.685 -0.18 0.925 0.32 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.07 1.315 7.67 1.315 7.67 2.17 6.26 2.17 6.26 1.89 6.56 1.89 6.56 2.05 7.55 2.05 7.55 0.62 7.42 0.62 7.42 0.48 6.26 0.48 6.26 0.36 7.54 0.36 7.54 0.5 7.67 0.5 7.67 1.195 7.83 1.195 7.83 1.075 8.07 1.075 ;
      POLYGON 7.43 0.86 7.345 0.86 7.345 1.81 7.43 1.81 7.43 1.93 7.19 1.93 7.19 1.81 7.225 1.81 7.225 0.86 7.19 0.86 7.19 0.74 7.43 0.74 ;
      POLYGON 7.05 1.77 7.04 1.77 7.04 1.79 6.8 1.79 6.8 1.77 4.275 1.77 4.275 1.65 5.095 1.65 5.095 0.72 4.525 0.72 4.525 0.6 5.215 0.6 5.215 1.65 6.93 1.65 6.93 0.72 6.8 0.72 6.8 0.6 7.05 0.6 ;
      POLYGON 5.96 0.705 5.9 0.705 5.9 0.72 5.48 0.72 5.48 1.405 5.96 1.405 5.96 1.525 5.36 1.525 5.36 0.6 5.72 0.6 5.72 0.585 5.96 0.585 ;
      RECT 2.985 1.89 5.96 2.01 ;
      RECT 2.405 0.36 5.64 0.48 ;
      RECT 2.405 2.13 5.64 2.25 ;
      POLYGON 4.97 1.04 4.17 1.04 4.17 1.285 4.05 1.285 4.05 0.92 4.97 0.92 ;
      POLYGON 4.075 0.72 3.93 0.72 3.93 1.77 1.725 1.77 1.725 2.17 0.985 2.17 0.985 1.81 0.325 1.81 0.325 1.93 0.205 1.93 0.205 1.69 0.505 1.69 0.505 0.92 0.205 0.92 0.205 0.44 1.605 0.44 1.605 0.32 1.725 0.32 1.725 0.56 0.325 0.56 0.325 0.8 0.625 0.8 0.625 1.69 1.105 1.69 1.105 2.05 1.605 2.05 1.605 1.65 3.81 1.65 3.81 0.6 4.075 0.6 ;
      POLYGON 3.69 1.08 3.57 1.08 3.57 1.02 2.81 1.02 2.81 1.16 2.885 1.16 2.885 1.28 2.645 1.28 2.645 1.16 2.69 1.16 2.69 0.9 3.57 0.9 3.57 0.84 3.69 0.84 ;
      POLYGON 3.225 1.53 1.94 1.53 1.94 0.6 3.205 0.6 3.205 0.72 2.06 0.72 2.06 1.41 3.225 1.41 ;
      POLYGON 1.485 1.52 1.405 1.52 1.405 1.81 1.465 1.81 1.465 1.93 1.225 1.93 1.225 1.81 1.285 1.81 1.285 1.52 1.245 1.52 1.245 1.4 1.285 1.4 1.285 0.8 1.225 0.8 1.225 0.68 1.465 0.68 1.465 0.8 1.405 0.8 1.405 1.4 1.485 1.4 ;
  END
END XNOR3X1

MACRO SEDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFXL 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.955 0.5 2.075 1.49 ;
        RECT 1.815 0.5 2.075 0.62 ;
        RECT 1.015 0.42 1.935 0.54 ;
        RECT 1.155 0.98 1.275 1.22 ;
        RECT 0.595 0.98 1.275 1.1 ;
        RECT 0.355 0.97 1.145 1.09 ;
        RECT 0.885 0.94 1.145 1.1 ;
        RECT 1.015 0.42 1.135 1.1 ;
        RECT 0.355 0.97 0.475 1.21 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.22 1.015 1.41 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.22 4.05 1.34 ;
        RECT 3.93 1.1 4.05 1.34 ;
        RECT 3.55 1.175 3.7 1.435 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 1.04 5.73 1.49 ;
        RECT 5.59 1.04 5.71 1.515 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.145 1.06 11.29 1.375 ;
        RECT 11.09 1.115 11.265 1.435 ;
    END
  END CK
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 1.59 2.98 1.83 ;
        RECT 2.71 1.59 2.98 1.71 ;
        RECT 2.71 0.885 2.83 1.71 ;
        RECT 2.68 0.885 2.83 1.145 ;
        RECT 2.535 0.885 2.83 1.005 ;
        RECT 2.535 0.6 2.655 1.005 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.19 1.69 6.45 1.81 ;
        RECT 6.16 1.465 6.31 1.725 ;
        RECT 6.19 0.8 6.31 1.81 ;
        RECT 6.09 0.68 6.21 0.92 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.01 -0.18 11.13 0.7 ;
        RECT 9.02 0.49 9.26 0.61 ;
        RECT 9.14 -0.18 9.26 0.61 ;
        RECT 7.2 0.49 7.44 0.61 ;
        RECT 7.32 -0.18 7.44 0.61 ;
        RECT 5.61 -0.18 5.73 0.92 ;
        RECT 3.73 -0.18 3.85 0.92 ;
        RECT 2.055 -0.18 2.175 0.38 ;
        RECT 0.615 -0.18 0.735 0.82 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 11.01 2 11.25 2.12 ;
        RECT 11.01 2 11.13 2.79 ;
        RECT 8.9 2.29 9.14 2.79 ;
        RECT 7.18 1.63 7.3 2.79 ;
        RECT 5.73 2.17 5.97 2.29 ;
        RECT 5.73 2.17 5.85 2.79 ;
        RECT 3.67 2.2 3.91 2.79 ;
        RECT 2.495 2.23 2.615 2.79 ;
        RECT 0.615 1.77 0.855 1.89 ;
        RECT 0.615 1.77 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.73 1.7 10.97 1.7 10.97 1.88 10.8 1.88 10.8 2.23 9.44 2.23 9.44 2.17 7.82 2.17 7.82 2.03 8.06 2.03 8.06 2.05 9.68 2.05 9.68 2.11 10.68 2.11 10.68 1.76 10.85 1.76 10.85 0.82 11.25 0.82 11.25 0.7 11.43 0.7 11.43 0.46 11.55 0.46 11.55 0.82 11.37 0.82 11.37 0.94 10.97 0.94 10.97 1.58 11.73 1.58 ;
      POLYGON 10.71 1.64 10.56 1.64 10.56 1.99 9.96 1.99 9.96 1.93 8.18 1.93 8.18 1.37 7.7 1.37 7.7 1.25 8.18 1.25 8.18 1.21 8.52 1.21 8.52 1.33 8.3 1.33 8.3 1.81 9.96 1.81 9.96 1.37 9.84 1.37 9.84 1.25 10.08 1.25 10.08 1.87 10.44 1.87 10.44 1.52 10.59 1.52 10.59 0.46 10.71 0.46 ;
      POLYGON 10.32 1.75 10.2 1.75 10.2 0.48 9.525 0.48 9.525 0.85 8.78 0.85 8.78 0.48 7.68 0.48 7.68 0.85 6.96 0.85 6.96 0.48 6.285 0.48 6.285 0.56 5.97 0.56 5.97 1.755 5.27 1.755 5.27 1.81 4.95 1.81 4.95 0.86 4.91 0.86 4.91 0.74 5.15 0.74 5.15 0.86 5.07 0.86 5.07 1.635 5.85 1.635 5.85 0.44 6.165 0.44 6.165 0.36 7.08 0.36 7.08 0.73 7.56 0.73 7.56 0.36 8.9 0.36 8.9 0.73 9.405 0.73 9.405 0.36 10.32 0.36 ;
      POLYGON 9.96 1.09 9.72 1.09 9.72 1.57 9.84 1.57 9.84 1.69 9.6 1.69 9.6 1.45 9.04 1.45 9.04 1.37 8.88 1.37 8.88 1.25 9.16 1.25 9.16 1.33 9.6 1.33 9.6 0.97 9.72 0.97 9.72 0.6 9.96 0.6 ;
      POLYGON 9.4 1.21 9.28 1.21 9.28 1.13 8.76 1.13 8.76 1.69 8.42 1.69 8.42 1.57 8.64 1.57 8.64 1.09 8.42 1.09 8.42 0.6 8.66 0.6 8.66 0.97 8.76 0.97 8.76 1.01 9.28 1.01 9.28 0.97 9.4 0.97 ;
      POLYGON 8.24 0.72 8.12 0.72 8.12 1.09 7.58 1.09 7.58 1.49 7.88 1.49 7.88 1.57 8 1.57 8 1.69 7.76 1.69 7.76 1.61 7.46 1.61 7.46 1.33 6.74 1.33 6.74 1.21 7.46 1.21 7.46 0.97 8 0.97 8 0.6 8.24 0.6 ;
      POLYGON 7.34 1.09 6.62 1.09 6.62 1.45 6.78 1.45 6.78 1.87 6.77 1.87 6.77 2.05 6.33 2.05 6.33 2.25 6.09 2.25 6.09 2.05 5.445 2.05 5.445 2.11 4.265 2.11 4.265 2.08 3.35 2.08 3.35 1.96 4.385 1.96 4.385 1.99 5.325 1.99 5.325 1.93 6.65 1.93 6.65 1.75 6.66 1.75 6.66 1.57 6.5 1.57 6.5 0.6 6.84 0.6 6.84 0.72 6.62 0.72 6.62 0.97 7.34 0.97 ;
      POLYGON 5.43 1.47 5.19 1.47 5.19 1.35 5.27 1.35 5.27 0.62 4.27 0.62 4.27 0.8 4.29 0.8 4.29 1.48 4.39 1.48 4.39 1.6 4.15 1.6 4.15 1.48 4.17 1.48 4.17 0.92 4.15 0.92 4.15 0.5 4.75 0.5 4.75 0.4 4.99 0.4 4.99 0.5 5.39 0.5 5.39 1.35 5.43 1.35 ;
      POLYGON 4.79 1.87 4.67 1.87 4.67 1.84 3.22 1.84 3.22 2.07 1.735 2.07 1.735 1.83 1.715 1.83 1.715 0.86 1.255 0.86 1.255 0.66 1.495 0.66 1.495 0.74 1.835 0.74 1.835 1.71 1.855 1.71 1.855 1.95 3.1 1.95 3.1 1.72 4.67 1.72 4.67 0.86 4.49 0.86 4.49 0.74 4.79 0.74 ;
      POLYGON 3.43 1.6 3.19 1.6 3.19 1.48 3.31 1.48 3.31 0.68 2.825 0.68 2.825 0.48 2.415 0.48 2.415 1.16 2.295 1.16 2.295 0.36 2.945 0.36 2.945 0.56 3.43 0.56 ;
      POLYGON 1.595 1.65 0.375 1.65 0.375 1.83 0.255 1.83 0.255 1.71 0.115 1.71 0.115 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.84 0.235 0.84 0.235 1.53 1.475 1.53 1.475 1.25 1.595 1.25 ;
  END
END SEDFFXL

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.955 1.24 2.075 1.48 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.84 1.36 2.075 1.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.71 1.575 0.83 ;
        RECT 1.395 1.32 1.515 2.21 ;
        RECT 0.515 0.76 1.455 0.88 ;
        RECT 0.515 1.32 1.515 1.44 ;
        RECT 0.555 1.32 0.8 1.725 ;
        RECT 0.555 1.32 0.675 2.21 ;
        RECT 0.555 0.64 0.675 0.88 ;
        RECT 0.515 0.76 0.635 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.815 -0.18 1.935 0.7 ;
        RECT 0.915 0.52 1.155 0.64 ;
        RECT 0.915 -0.18 1.035 0.64 ;
        RECT 0.135 -0.18 0.255 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.815 1.845 1.935 2.79 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.355 2.21 2.235 2.21 2.235 1.12 1.415 1.12 1.415 1.17 1.175 1.17 1.175 1.12 0.995 1.12 0.995 1.17 0.755 1.17 0.755 1.05 0.875 1.05 0.875 1 2.235 1 2.235 0.65 2.355 0.65 ;
  END
END BUFX4

MACRO AOI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X1 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.095 1.67 1.435 ;
        RECT 1.48 0.975 1.6 1.315 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.01 1.18 1.15 ;
        RECT 0.94 1.01 1.09 1.435 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.98 0.8 1.435 ;
        RECT 0.68 0.96 0.8 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.78 0.51 1.15 ;
        RECT 0.32 0.815 0.44 1.19 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.44 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 1.555 1.91 1.675 ;
        RECT 1.79 0.72 1.91 1.675 ;
        RECT 0.86 0.72 1.91 0.84 ;
        RECT 1.64 1.555 1.76 2.21 ;
        RECT 1.52 0.6 1.76 0.84 ;
        RECT 1.52 0.595 1.67 0.855 ;
        RECT 0.74 0.67 0.98 0.79 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 1.16 0.48 1.4 0.6 ;
        RECT 1.16 -0.18 1.28 0.6 ;
        RECT 0.16 -0.18 0.28 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 0.58 1.795 0.7 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.12 2.21 1 2.21 1 1.675 0.28 1.675 0.28 2.21 0.16 2.21 0.16 1.555 1.12 1.555 ;
  END
END AOI211X1

MACRO TLATX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX4 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.045 0.51 1.44 ;
        RECT 0.39 0.835 0.51 1.44 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 1.46 8.63 1.775 ;
        RECT 8.325 1.46 8.63 1.77 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.125 1.32 2.245 2.21 ;
        RECT 1.26 1.32 2.245 1.44 ;
        RECT 1.025 0.8 2.105 0.92 ;
        RECT 1.985 0.68 2.105 0.92 ;
        RECT 1.285 0.8 1.405 2.21 ;
        RECT 1.23 1.175 1.405 1.435 ;
        RECT 1.025 0.68 1.145 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.825 0.8 5.945 0.92 ;
        RECT 5.825 0.68 5.945 0.92 ;
        RECT 5.485 1.32 5.605 2.21 ;
        RECT 4.71 1.32 5.605 1.44 ;
        RECT 4.865 0.68 4.985 0.92 ;
        RECT 4.71 1.175 4.945 1.56 ;
        RECT 4.825 0.8 4.945 1.56 ;
        RECT 4.645 1.44 4.765 2.21 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 8.545 -0.18 8.665 0.38 ;
        RECT 7.265 -0.18 7.385 0.4 ;
        RECT 6.245 -0.18 6.485 0.32 ;
        RECT 5.285 -0.18 5.525 0.32 ;
        RECT 4.325 -0.18 4.565 0.32 ;
        RECT 3.365 -0.18 3.605 0.32 ;
        RECT 2.405 -0.18 2.645 0.32 ;
        RECT 1.445 -0.18 1.685 0.32 ;
        RECT 0.545 -0.18 0.665 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 8.385 1.92 8.505 2.79 ;
        RECT 6.805 1.82 6.925 2.79 ;
        RECT 5.905 1.56 6.025 2.79 ;
        RECT 5.065 1.56 5.185 2.79 ;
        RECT 4.225 1.56 4.345 2.79 ;
        RECT 3.385 1.56 3.505 2.79 ;
        RECT 2.545 1.56 2.665 2.79 ;
        RECT 1.705 1.56 1.825 2.79 ;
        RECT 0.865 1.56 0.985 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.205 0.86 9.085 0.86 9.085 1.34 8.925 1.34 8.925 2.04 8.805 2.04 8.805 1.34 8.125 1.34 8.125 1.58 7.585 1.58 7.585 1.7 7.465 1.7 7.465 1.46 8.005 1.46 8.005 1.22 8.965 1.22 8.965 0.74 9.205 0.74 ;
      POLYGON 9.045 0.52 8.925 0.52 8.925 0.62 7.645 0.62 7.645 0.64 7.025 0.64 7.025 0.56 0.905 0.56 0.905 0.68 0.255 0.68 0.255 0.92 0.24 0.92 0.24 1.56 0.505 1.56 0.505 1.8 0.385 1.8 0.385 1.68 0.12 1.68 0.12 0.8 0.135 0.8 0.135 0.56 0.785 0.56 0.785 0.44 7.145 0.44 7.145 0.52 7.525 0.52 7.525 0.5 7.645 0.5 7.645 0.42 7.885 0.42 7.885 0.5 8.805 0.5 8.805 0.4 9.045 0.4 ;
      POLYGON 8.025 0.86 7.885 0.86 7.885 1.34 7.345 1.34 7.345 1.82 7.585 1.82 7.585 1.86 7.705 1.86 7.705 1.98 7.465 1.98 7.465 1.94 7.225 1.94 7.225 1.7 6.625 1.7 6.625 1.37 6.745 1.37 6.745 1.58 7.225 1.58 7.225 1.22 7.765 1.22 7.765 0.74 8.025 0.74 ;
      POLYGON 7.105 1.46 6.985 1.46 6.985 1.25 6.785 1.25 6.785 1.2 6.505 1.2 6.505 2.21 6.385 2.21 6.385 1.2 5.625 1.2 5.625 1.08 6.785 1.08 6.785 0.68 6.905 0.68 6.905 1.13 7.105 1.13 ;
      POLYGON 4.025 0.92 3.065 0.92 3.065 1.08 3.085 1.08 3.085 1.32 3.925 1.32 3.925 2.21 3.805 2.21 3.805 1.44 3.085 1.44 3.085 2.21 2.965 2.21 2.965 1.2 1.925 1.2 1.925 1.08 2.945 1.08 2.945 0.68 3.065 0.68 3.065 0.8 3.905 0.8 3.905 0.68 4.025 0.68 ;
  END
END TLATX4

MACRO BUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX20 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.54 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.02 1.26 8.62 1.38 ;
        RECT 8.135 1.23 8.395 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6387 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.96 1.425 7.08 2.21 ;
        RECT 0.36 0.945 7.08 1.065 ;
        RECT 6.96 0.4 7.08 1.065 ;
        RECT 0.24 1.425 7.08 1.545 ;
        RECT 6.12 1.425 6.24 2.21 ;
        RECT 6.12 0.4 6.24 1.065 ;
        RECT 5.28 1.425 5.4 2.21 ;
        RECT 5.22 0.4 5.34 1.065 ;
        RECT 4.44 1.425 4.56 2.21 ;
        RECT 4.38 0.4 4.5 1.065 ;
        RECT 3.6 1.425 3.72 2.21 ;
        RECT 3.54 0.4 3.66 1.065 ;
        RECT 2.76 1.425 2.88 2.21 ;
        RECT 2.7 0.4 2.82 1.065 ;
        RECT 1.92 1.425 2.04 2.21 ;
        RECT 1.86 0.4 1.98 1.065 ;
        RECT 1.08 1.425 1.2 2.21 ;
        RECT 1.02 0.4 1.14 1.065 ;
        RECT 0.36 0.945 0.51 1.545 ;
        RECT 0.36 0.785 0.48 1.545 ;
        RECT 0.24 1.425 0.36 2.21 ;
        RECT 0.18 0.785 0.48 0.905 ;
        RECT 0.18 0.4 0.3 0.905 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.06 -0.18 9.18 0.72 ;
        RECT 8.22 -0.18 8.34 0.72 ;
        RECT 7.38 -0.18 7.5 0.91 ;
        RECT 6.54 -0.18 6.66 0.825 ;
        RECT 5.64 -0.18 5.76 0.825 ;
        RECT 4.8 -0.18 4.92 0.825 ;
        RECT 3.96 -0.18 4.08 0.825 ;
        RECT 3.12 -0.18 3.24 0.825 ;
        RECT 2.28 -0.18 2.4 0.825 ;
        RECT 1.44 -0.18 1.56 0.825 ;
        RECT 0.6 -0.18 0.72 0.825 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.06 1.74 9.18 2.79 ;
        RECT 8.22 1.74 8.34 2.79 ;
        RECT 7.38 1.56 7.5 2.79 ;
        RECT 6.54 1.665 6.66 2.79 ;
        RECT 5.7 1.665 5.82 2.79 ;
        RECT 4.86 1.665 4.98 2.79 ;
        RECT 4.02 1.665 4.14 2.79 ;
        RECT 3.18 1.665 3.3 2.79 ;
        RECT 2.34 1.665 2.46 2.79 ;
        RECT 1.5 1.665 1.62 2.79 ;
        RECT 0.66 1.665 0.78 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.6 0.96 7.9 0.96 7.9 1.5 9.6 1.5 9.6 2.21 9.48 2.21 9.48 1.62 8.76 1.62 8.76 2.21 8.64 2.21 8.64 1.62 7.92 1.62 7.92 2.21 7.8 2.21 7.8 1.62 7.78 1.62 7.78 1.305 0.82 1.305 0.82 1.185 7.78 1.185 7.78 0.84 7.8 0.84 7.8 0.67 7.92 0.67 7.92 0.84 8.64 0.84 8.64 0.67 8.76 0.67 8.76 0.84 9.48 0.84 9.48 0.67 9.6 0.67 ;
  END
END BUFX20

MACRO NAND2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.76 0.51 1.24 ;
        RECT 0.36 0.76 0.51 1.215 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1 1.38 1.5 ;
        RECT 1.23 1 1.38 1.47 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3284 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.62 1.36 0.74 2.21 ;
        RECT 0.12 1.36 0.74 1.48 ;
        RECT 0.12 0.52 0.46 0.64 ;
        RECT 0.34 0.4 0.46 0.64 ;
        RECT 0.07 1.175 0.24 1.435 ;
        RECT 0.12 0.52 0.24 1.48 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.98 -0.18 1.1 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.04 1.62 1.16 2.79 ;
        RECT 0.2 1.6 0.32 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.62 1.74 1.58 1.74 1.58 1.86 1.46 1.86 1.46 1.62 1.5 1.62 1.5 0.88 1.11 0.88 1.11 1.09 0.84 1.09 0.84 0.97 0.99 0.97 0.99 0.76 1.46 0.76 1.46 0.59 1.58 0.59 1.58 0.71 1.62 0.71 ;
  END
END NAND2BX1

MACRO OAI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211XL 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.31 1.25 1.48 1.49 ;
        RECT 1.23 1.175 1.43 1.435 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 1.17 1.11 1.595 ;
        RECT 0.94 1.17 1.11 1.58 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.8 1.63 ;
        RECT 0.67 1.17 0.79 1.65 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.465 0.51 1.865 ;
        RECT 0.35 1.17 0.47 1.585 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 1.71 1.895 1.95 ;
        RECT 1.615 0.57 1.735 0.81 ;
        RECT 1.6 0.69 1.72 1.95 ;
        RECT 1.52 1.755 1.67 2.015 ;
        RECT 0.77 1.77 1.895 1.89 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 0.555 -0.18 0.675 0.81 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.31 2.23 1.43 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.155 0.75 1.035 0.75 1.035 1.05 0.195 1.05 0.195 0.75 0.075 0.75 0.075 0.63 0.315 0.63 0.315 0.93 0.915 0.93 0.915 0.63 1.155 0.63 ;
  END
END OAI211XL

MACRO OA22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X1 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.255 1.295 ;
        RECT 1.135 1.055 1.255 1.295 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.165 0.51 1.62 ;
        RECT 0.38 1.1 0.5 1.62 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1 0.82 1.435 ;
        RECT 0.7 0.98 0.82 1.435 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.615 1.4 1.93 1.52 ;
        RECT 1.615 1.28 1.735 1.52 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.42 0.65 2.825 0.77 ;
        RECT 2.42 0.65 2.54 1.145 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.275 1.005 2.395 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 2.165 -0.18 2.285 0.53 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.855 1.845 1.975 2.79 ;
        RECT 0.22 1.74 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.155 1.18 1.855 1.18 1.855 1.16 1.495 1.16 1.495 1.8 0.995 1.8 0.995 1.68 1.375 1.68 1.375 0.8 1.475 0.8 1.475 0.68 1.595 0.68 1.595 0.92 1.495 0.92 1.495 1.04 1.975 1.04 1.975 1.06 2.155 1.06 ;
      POLYGON 2.015 0.92 1.895 0.92 1.895 0.56 1.175 0.56 1.175 0.92 1.055 0.92 1.055 0.86 0.075 0.86 0.075 0.74 1.055 0.74 1.055 0.44 2.015 0.44 ;
  END
END OA22X1

MACRO CLKINVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX4 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 1.26 1.4 1.38 ;
        RECT 0.885 1.23 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.52 0.85 1.64 1.725 ;
        RECT 1.5 1.5 1.62 2.21 ;
        RECT 0.66 0.85 1.64 0.97 ;
        RECT 1.5 0.68 1.62 0.97 ;
        RECT 0.66 1.5 1.67 1.62 ;
        RECT 0.66 1.5 0.78 2.21 ;
        RECT 0.66 0.68 0.78 0.97 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.92 -0.18 2.04 0.73 ;
        RECT 1.08 -0.18 1.2 0.73 ;
        RECT 0.24 -0.18 0.36 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.92 1.56 2.04 2.79 ;
        RECT 1.08 1.74 1.2 2.79 ;
        RECT 0.24 1.56 0.36 2.79 ;
    END
  END VDD
END CLKINVX4

MACRO AOI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X4 0 0 ;
  SIZE 10.73 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.855 0.75 9.975 1.17 ;
        RECT 5.375 0.75 9.975 0.87 ;
        RECT 7.5 0.75 7.74 1.09 ;
        RECT 5.235 0.94 5.495 1.09 ;
        RECT 5.375 0.75 5.495 1.09 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.755 0.75 4.875 1.15 ;
        RECT 4.71 0.75 4.875 1.145 ;
        RECT 0.575 0.75 4.875 0.87 ;
        RECT 2.64 0.75 2.88 1.09 ;
        RECT 0.575 0.75 0.695 1.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.29 0.99 4.59 1.11 ;
        RECT 2.4 1.21 3.435 1.33 ;
        RECT 3.29 0.99 3.435 1.33 ;
        RECT 2.4 1.06 2.52 1.33 ;
        RECT 1.34 1.06 2.52 1.18 ;
        RECT 0.855 1.175 1.46 1.295 ;
        RECT 1.23 1.175 1.38 1.435 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.35 1.175 9.655 1.38 ;
        RECT 9.535 1.14 9.655 1.38 ;
        RECT 9.35 1.175 9.5 1.435 ;
        RECT 9.01 1.175 9.655 1.295 ;
        RECT 9.01 1.04 9.13 1.295 ;
        RECT 7.86 1.04 9.13 1.16 ;
        RECT 7.065 1.21 7.98 1.33 ;
        RECT 7.86 1.04 7.98 1.33 ;
        RECT 7.065 0.99 7.185 1.33 ;
        RECT 5.795 0.99 7.185 1.11 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.635 1.28 8.875 1.4 ;
        RECT 6.78 1.45 8.755 1.57 ;
        RECT 8.635 1.28 8.755 1.57 ;
        RECT 6.78 1.23 6.945 1.57 ;
        RECT 6.635 1.28 6.945 1.4 ;
        RECT 6.685 1.23 6.945 1.4 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.23 4.045 1.38 ;
        RECT 2.16 1.45 3.87 1.57 ;
        RECT 3.75 1.26 3.905 1.48 ;
        RECT 2.16 1.3 2.28 1.57 ;
        RECT 1.615 1.3 2.28 1.42 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.7984 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.795 1.56 9.915 2.01 ;
        RECT 5.595 1.69 9.915 1.81 ;
        RECT 8.955 1.56 9.075 2.01 ;
        RECT 1.535 0.51 8.935 0.63 ;
        RECT 8.115 1.69 8.235 2.01 ;
        RECT 7.275 1.69 7.395 2.01 ;
        RECT 6.435 1.56 6.555 2.01 ;
        RECT 5.595 1.23 5.715 2.01 ;
        RECT 4.995 1.23 5.715 1.38 ;
        RECT 4.995 1.18 5.15 1.43 ;
        RECT 4.995 0.51 5.115 1.43 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.73 0.18 ;
        RECT 9.955 0.46 10.195 0.58 ;
        RECT 9.955 -0.18 10.075 0.58 ;
        RECT 7.675 -0.18 7.915 0.39 ;
        RECT 5.035 -0.18 5.275 0.39 ;
        RECT 2.555 -0.18 2.795 0.39 ;
        RECT 0.375 0.46 0.615 0.58 ;
        RECT 0.375 -0.18 0.495 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.73 2.79 ;
        RECT 4.755 1.93 4.875 2.79 ;
        RECT 3.915 1.93 4.035 2.79 ;
        RECT 3.075 1.93 3.195 2.79 ;
        RECT 2.235 1.93 2.355 2.79 ;
        RECT 1.395 1.93 1.515 2.79 ;
        RECT 0.555 1.93 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.335 2.25 5.175 2.25 5.175 1.81 4.455 1.81 4.455 2.21 4.335 2.21 4.335 1.81 3.615 1.81 3.615 2.21 3.495 2.21 3.495 1.81 2.775 1.81 2.775 2.21 2.655 2.21 2.655 1.81 1.935 1.81 1.935 2.21 1.815 2.21 1.815 1.81 1.095 1.81 1.095 2.21 0.975 2.21 0.975 1.81 0.255 1.81 0.255 2.21 0.135 2.21 0.135 1.56 0.255 1.56 0.255 1.69 0.975 1.69 0.975 1.56 1.095 1.56 1.095 1.69 1.815 1.69 1.815 1.56 1.935 1.56 1.935 1.69 4.335 1.69 4.335 1.56 4.455 1.56 4.455 1.69 5.175 1.69 5.175 1.56 5.295 1.56 5.295 2.13 6.015 2.13 6.015 1.93 6.135 1.93 6.135 2.13 6.855 2.13 6.855 1.93 6.975 1.93 6.975 2.13 7.695 2.13 7.695 1.93 7.815 1.93 7.815 2.13 8.535 2.13 8.535 1.93 8.655 1.93 8.655 2.13 9.375 2.13 9.375 1.93 9.495 1.93 9.495 2.13 10.215 2.13 10.215 1.56 10.335 1.56 ;
  END
END AOI33X4

MACRO TBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX16 0 0 ;
  SIZE 16.53 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2184 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.54 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.4044 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 0.85 1.635 1.1 ;
        RECT 0.555 0.85 1.635 0.97 ;
        RECT 0.36 0.885 0.675 1.125 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.855 1.185 9.095 1.305 ;
        RECT 8.855 1 8.975 1.305 ;
        RECT 5.515 1 8.975 1.12 ;
        RECT 5.515 0.76 5.635 1.12 ;
        RECT 4.935 0.76 5.635 0.88 ;
        RECT 4.935 0.41 5.055 0.88 ;
        RECT 4.335 0.41 5.055 0.53 ;
        RECT 3.855 0.795 4.455 0.915 ;
        RECT 4.335 0.41 4.455 0.915 ;
        RECT 4.12 0.795 4.24 1.15 ;
        RECT 3.855 0.36 3.975 0.915 ;
        RECT 3.155 0.36 3.975 0.48 ;
        RECT 2.45 0.71 3.275 0.83 ;
        RECT 3.155 0.36 3.275 0.83 ;
        RECT 2.715 0.71 2.835 1.12 ;
        RECT 2.45 0.36 2.57 0.83 ;
        RECT 1.755 0.36 2.57 0.48 ;
        RECT 1.755 0.94 2.015 1.09 ;
        RECT 1.175 1.22 1.875 1.34 ;
        RECT 1.755 0.36 1.875 1.34 ;
        RECT 0.795 1.15 1.295 1.27 ;
        RECT 1.175 1.09 1.295 1.34 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.7648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.695 1.32 15.815 2.21 ;
        RECT 15.675 0.59 15.795 1.44 ;
        RECT 9.93 1.32 15.815 1.44 ;
        RECT 13.995 0.76 15.795 0.88 ;
        RECT 14.855 1.32 14.975 2.21 ;
        RECT 14.835 0.59 14.955 0.88 ;
        RECT 14.015 1.32 14.135 2.21 ;
        RECT 13.995 0.59 14.115 0.88 ;
        RECT 13.175 1.32 13.295 2.21 ;
        RECT 13.155 0.59 13.275 1.44 ;
        RECT 12.315 0.76 13.275 0.88 ;
        RECT 12.335 1.32 12.455 2.21 ;
        RECT 12.315 0.59 12.435 0.88 ;
        RECT 11.495 1.32 11.615 2.21 ;
        RECT 11.475 0.59 11.595 0.83 ;
        RECT 11.295 0.71 11.595 0.83 ;
        RECT 11.295 0.71 11.415 1.44 ;
        RECT 10.635 0.76 11.415 0.88 ;
        RECT 10.655 1.32 10.775 2.21 ;
        RECT 10.635 0.59 10.755 0.88 ;
        RECT 9.93 1.175 10.08 1.44 ;
        RECT 9.93 0.96 10.05 1.68 ;
        RECT 9.815 1.56 9.935 2.21 ;
        RECT 9.795 0.96 10.05 1.08 ;
        RECT 9.795 0.59 9.915 1.08 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 16.53 0.18 ;
        RECT 16.095 -0.18 16.215 0.64 ;
        RECT 15.255 -0.18 15.375 0.64 ;
        RECT 14.415 -0.18 14.535 0.64 ;
        RECT 13.575 -0.18 13.695 0.64 ;
        RECT 12.735 -0.18 12.855 0.64 ;
        RECT 11.895 -0.18 12.015 0.64 ;
        RECT 11.055 -0.18 11.175 0.64 ;
        RECT 10.215 -0.18 10.335 0.64 ;
        RECT 9.375 -0.18 9.495 0.64 ;
        RECT 8.535 -0.18 8.655 0.64 ;
        RECT 7.695 -0.18 7.815 0.64 ;
        RECT 6.855 -0.18 6.975 0.64 ;
        RECT 6.015 -0.18 6.135 0.64 ;
        RECT 5.175 -0.18 5.295 0.64 ;
        RECT 4.095 -0.18 4.215 0.675 ;
        RECT 2.695 0.47 2.935 0.59 ;
        RECT 2.695 -0.18 2.815 0.59 ;
        RECT 0.955 -0.18 1.075 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 16.53 2.79 ;
        RECT 16.115 1.56 16.235 2.79 ;
        RECT 15.275 1.56 15.395 2.79 ;
        RECT 14.435 1.56 14.555 2.79 ;
        RECT 13.595 1.56 13.715 2.79 ;
        RECT 12.755 1.56 12.875 2.79 ;
        RECT 11.915 1.56 12.035 2.79 ;
        RECT 11.075 1.56 11.195 2.79 ;
        RECT 10.235 1.56 10.355 2.79 ;
        RECT 8.995 1.96 9.235 2.08 ;
        RECT 8.995 1.96 9.115 2.79 ;
        RECT 7.715 1.96 7.955 2.08 ;
        RECT 7.715 1.96 7.835 2.79 ;
        RECT 6.435 1.96 6.675 2.08 ;
        RECT 6.435 1.96 6.555 2.79 ;
        RECT 4.735 1.53 4.855 2.79 ;
        RECT 4.615 1.53 4.855 1.93 ;
        RECT 3.835 1.72 3.955 2.79 ;
        RECT 2.935 2.23 3.055 2.79 ;
        RECT 2.035 1.72 2.155 2.79 ;
        RECT 1.135 2.23 1.255 2.79 ;
        RECT 0.235 1.72 0.355 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.795 1.44 9.695 1.44 9.695 1.84 8.775 1.84 8.775 2.25 8.075 2.25 8.075 1.84 7.545 1.84 7.545 2.25 6.895 2.25 6.895 1.84 6.275 1.84 6.275 2.25 4.975 2.25 4.975 1.41 4.375 1.41 4.375 1.99 4.255 1.99 4.255 1.6 3.535 1.6 3.535 1.95 3.415 1.95 3.415 1.6 2.575 1.6 2.575 1.98 2.455 1.98 2.455 1.6 1.735 1.6 1.735 1.95 1.615 1.95 1.615 1.6 0.775 1.6 0.775 2.21 0.655 2.21 0.655 1.6 0.12 1.6 0.12 0.645 0.315 0.645 0.315 0.525 0.435 0.525 0.435 0.765 0.24 0.765 0.24 1.48 1.615 1.48 1.615 1.46 1.735 1.46 1.735 1.48 2.135 1.48 2.135 0.72 1.995 0.72 1.995 0.6 2.255 0.6 2.255 1.48 3.615 1.48 3.615 0.72 3.395 0.72 3.395 0.6 3.735 0.6 3.735 1.48 4.255 1.48 4.255 1.29 5.095 1.29 5.095 2.13 6.155 2.13 6.155 1.72 7.015 1.72 7.015 2.13 7.425 2.13 7.425 1.72 8.195 1.72 8.195 2.13 8.655 2.13 8.655 1.72 9.575 1.72 9.575 1.32 9.675 1.32 9.675 1.2 9.795 1.2 ;
      POLYGON 9.455 1.225 9.335 1.225 9.335 1.6 8.535 1.6 8.535 2.01 8.415 2.01 8.415 1.6 7.255 1.6 7.255 2.01 7.135 2.01 7.135 1.6 6.035 1.6 6.035 2.01 5.795 2.01 5.795 1.68 5.915 1.68 5.915 1.48 9.215 1.48 9.215 0.88 5.755 0.88 5.755 0.64 5.595 0.64 5.595 0.4 5.715 0.4 5.715 0.52 5.875 0.52 5.875 0.76 6.435 0.76 6.435 0.505 6.555 0.505 6.555 0.76 7.275 0.76 7.275 0.505 7.395 0.505 7.395 0.76 8.115 0.76 8.115 0.505 8.235 0.505 8.235 0.76 8.955 0.76 8.955 0.505 9.075 0.505 9.075 0.76 9.335 0.76 9.335 1.105 9.455 1.105 ;
      POLYGON 8.455 1.36 5.515 1.36 5.515 1.93 5.275 1.93 5.275 1.12 4.575 1.12 4.575 0.65 4.815 0.65 4.815 1 5.395 1 5.395 1.24 8.455 1.24 ;
      POLYGON 3.495 1.36 2.375 1.36 2.375 1.12 2.495 1.12 2.495 1.24 3.255 1.24 3.255 0.95 3.495 0.95 ;
  END
END TBUFX16

MACRO SDFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX1 0 0 ;
  SIZE 10.73 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.845 1.34 2.125 1.46 ;
        RECT 2.005 1.22 2.125 1.46 ;
        RECT 1.81 1.465 1.965 1.725 ;
        RECT 1.845 1.34 1.965 1.725 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3456 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.88 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 1.205 3.525 1.425 ;
        RECT 3.205 1.205 3.465 1.45 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.19 0.76 8.445 0.96 ;
        RECT 8.19 0.76 8.34 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.585 0.94 9.845 1.17 ;
        RECT 9.665 0.94 9.785 1.35 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.005 0.885 10.37 1.145 ;
        RECT 10.005 0.7 10.125 1.145 ;
        RECT 9.345 0.7 10.125 0.82 ;
        RECT 8.805 1.03 9.465 1.15 ;
        RECT 9.345 0.7 9.465 1.15 ;
        RECT 8.805 1.03 8.925 1.27 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 2.21 ;
        RECT 1.23 0.885 1.485 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.73 0.18 ;
        RECT 9.765 0.46 10.005 0.58 ;
        RECT 9.765 -0.18 9.885 0.58 ;
        RECT 8.325 -0.18 8.445 0.64 ;
        RECT 5.765 0.47 6.005 0.59 ;
        RECT 5.885 -0.18 6.005 0.59 ;
        RECT 3.545 -0.18 3.665 0.605 ;
        RECT 1.725 0.55 1.965 0.67 ;
        RECT 1.725 -0.18 1.845 0.67 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.73 2.79 ;
        RECT 9.725 1.71 9.845 2.79 ;
        RECT 8.485 2.23 8.605 2.79 ;
        RECT 6.445 2.05 6.685 2.17 ;
        RECT 6.445 2.05 6.565 2.79 ;
        RECT 5.485 2.29 5.725 2.79 ;
        RECT 3.485 2.29 3.725 2.79 ;
        RECT 2.655 2.15 2.775 2.79 ;
        RECT 1.785 1.845 1.905 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.61 1.71 10.265 1.71 10.265 1.83 10.145 1.83 10.145 1.59 9.285 1.59 9.285 1.45 9.165 1.45 9.165 1.33 9.405 1.33 9.405 1.47 10.49 1.47 10.49 0.765 10.245 0.765 10.245 0.4 10.365 0.4 10.365 0.645 10.61 0.645 ;
      POLYGON 9.365 0.58 9.225 0.58 9.225 0.91 8.685 0.91 8.685 1.77 9.245 1.77 9.245 1.89 8.685 1.89 8.685 2.01 7.615 2.01 7.615 1.34 7.405 1.34 7.405 0.86 7.305 0.86 7.305 0.62 7.425 0.62 7.425 0.74 7.525 0.74 7.525 1.22 7.735 1.22 7.735 1.89 8.565 1.89 8.565 0.79 9.105 0.79 9.105 0.46 9.365 0.46 ;
      POLYGON 8.345 2.25 7.22 2.25 7.22 1.94 7.075 1.94 7.075 2.04 6.955 2.04 6.955 1.93 2.265 1.93 2.265 1.57 2.325 1.57 2.325 0.74 2.565 0.74 2.565 0.86 2.445 0.86 2.445 1.69 2.385 1.69 2.385 1.81 4.105 1.81 4.105 0.94 4.225 0.94 4.225 1.81 4.765 1.81 4.765 1.37 4.625 1.37 4.625 1.25 4.885 1.25 4.885 1.81 6.955 1.81 6.955 1.8 7.075 1.8 7.075 1.82 7.34 1.82 7.34 2.13 8.345 2.13 ;
      POLYGON 8.185 1.77 7.945 1.77 7.945 0.98 7.765 0.98 7.765 1.1 7.645 1.1 7.645 0.5 6.245 0.5 6.245 0.83 5.525 0.83 5.525 0.5 5.165 0.5 5.165 1.18 5.045 1.18 5.045 0.38 5.645 0.38 5.645 0.71 6.125 0.71 6.125 0.38 6.545 0.38 6.545 0.36 6.785 0.36 6.785 0.38 7.765 0.38 7.765 0.4 7.885 0.4 7.885 0.86 8.065 0.86 8.065 1.65 8.185 1.65 ;
      POLYGON 7.315 1.7 7.195 1.7 7.195 1.58 7.165 1.58 7.165 1.4 5.645 1.4 5.645 1.43 5.525 1.43 5.525 1.19 5.645 1.19 5.645 1.28 6.885 1.28 6.885 0.62 7.005 0.62 7.005 1.28 7.285 1.28 7.285 1.46 7.315 1.46 ;
      POLYGON 6.955 1.64 6.205 1.64 6.205 1.69 5.965 1.69 5.965 1.57 6.085 1.57 6.085 1.52 6.955 1.52 ;
      POLYGON 6.565 1.12 6.325 1.12 6.325 1.07 5.405 1.07 5.405 1.69 5.005 1.69 5.005 1.57 5.285 1.57 5.285 0.62 5.405 0.62 5.405 0.95 6.445 0.95 6.445 1 6.565 1 ;
      RECT 3.165 2.05 6.045 2.17 ;
      POLYGON 4.645 1.69 4.385 1.69 4.385 0.82 3.975 0.82 3.975 0.845 3.085 0.845 3.085 0.48 2.925 0.48 2.925 0.36 3.205 0.36 3.205 0.725 3.855 0.725 3.855 0.7 4.385 0.7 4.385 0.62 4.505 0.62 4.505 1.57 4.645 1.57 ;
      POLYGON 3.885 1.205 3.765 1.205 3.765 1.085 3.085 1.085 3.085 1.57 3.245 1.57 3.245 1.69 2.965 1.69 2.965 1.085 2.845 1.085 2.845 0.74 2.685 0.74 2.685 0.62 2.205 0.62 2.205 1.1 1.725 1.1 1.725 1.24 1.605 1.24 1.605 0.98 2.085 0.98 2.085 0.5 2.805 0.5 2.805 0.62 2.965 0.62 2.965 0.965 3.885 0.965 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END SDFFRX1

MACRO DFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX8 0 0 ;
  SIZE 13.63 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.465 2.775 2.21 ;
        RECT 2.655 0.68 2.775 1.005 ;
        RECT 2.635 0.885 2.755 1.585 ;
        RECT 0.07 1.005 2.755 1.125 ;
        RECT 1.815 0.68 1.935 2.21 ;
        RECT 0.975 0.68 1.095 2.205 ;
        RECT 0.135 0.68 0.255 2.205 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.02 5.15 1.435 ;
        RECT 5 0.92 5.12 1.435 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.32 2.13 9.825 2.25 ;
        RECT 9.32 1.76 9.44 2.25 ;
        RECT 8.565 1.76 9.44 1.88 ;
        RECT 7.085 2.13 8.685 2.25 ;
        RECT 8.565 1.76 8.685 2.25 ;
        RECT 7.085 1.76 7.205 2.25 ;
        RECT 6.235 1.76 7.205 1.88 ;
        RECT 5.705 1.89 6.355 2.01 ;
        RECT 6.235 1.76 6.355 2.01 ;
        RECT 5.705 1.23 5.825 2.01 ;
        RECT 5.58 1.175 5.73 1.435 ;
        RECT 5.61 1.11 5.73 1.435 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.905 0.895 12.165 1.13 ;
        RECT 11.825 1.01 12.065 1.22 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.12 1.16 13.27 1.58 ;
        RECT 13.125 1.04 13.245 1.58 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.63 0.18 ;
        RECT 13.375 -0.18 13.495 0.4 ;
        RECT 12.045 -0.18 12.285 0.32 ;
        RECT 10.505 -0.18 10.625 0.68 ;
        RECT 5.205 -0.18 5.445 0.32 ;
        RECT 3.915 -0.18 4.035 0.69 ;
        RECT 3.075 -0.18 3.195 0.69 ;
        RECT 2.235 -0.18 2.355 0.67 ;
        RECT 1.395 -0.18 1.515 0.67 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.63 2.79 ;
        RECT 13.3 1.7 13.42 2.79 ;
        RECT 12.025 1.58 12.145 2.79 ;
        RECT 10.52 1.86 10.64 2.79 ;
        RECT 10.4 1.86 10.64 2 ;
        RECT 8.925 2 9.045 2.79 ;
        RECT 8.805 2 9.045 2.12 ;
        RECT 6.725 2 6.965 2.12 ;
        RECT 6.725 2 6.845 2.79 ;
        RECT 5.225 1.795 5.345 2.79 ;
        RECT 5.105 1.795 5.345 1.915 ;
        RECT 3.915 1.56 4.035 2.79 ;
        RECT 3.075 1.56 3.195 2.79 ;
        RECT 2.235 1.465 2.355 2.79 ;
        RECT 1.395 1.465 1.515 2.79 ;
        RECT 0.555 1.465 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.095 0.92 13.005 0.92 13.005 1.04 13 1.04 13 1.82 12.88 1.82 12.88 0.92 12.885 0.92 12.885 0.8 12.975 0.8 12.975 0.56 11.705 0.56 11.705 1.12 11.565 1.12 11.565 0.88 11.585 0.88 11.585 0.48 11.065 0.48 11.065 1.14 11.185 1.14 11.185 1.26 10.945 1.26 10.945 0.92 9.645 0.92 9.645 1.16 8.405 1.16 8.405 1.04 9.525 1.04 9.525 0.8 10.945 0.8 10.945 0.36 11.705 0.36 11.705 0.44 12.405 0.44 12.405 0.36 12.645 0.36 12.645 0.44 13.095 0.44 ;
      POLYGON 12.765 0.8 12.645 0.8 12.645 1.46 12.565 1.46 12.565 1.82 12.445 1.82 12.445 1.46 11.665 1.46 11.665 2.25 10.76 2.25 10.76 1.74 10.28 1.74 10.28 2.01 9.56 2.01 9.56 1.64 8.445 1.64 8.445 2.01 7.365 2.01 7.365 1.08 7.485 1.08 7.485 1.89 7.845 1.89 7.845 0.96 7.925 0.96 7.925 0.84 8.045 0.84 8.045 1.08 7.965 1.08 7.965 1.89 8.325 1.89 8.325 1.52 9.68 1.52 9.68 1.89 10.16 1.89 10.16 1.62 10.88 1.62 10.88 2.13 11.545 2.13 11.545 1.24 11.665 1.24 11.665 1.34 12.525 1.34 12.525 0.68 12.765 0.68 ;
      POLYGON 11.465 0.72 11.425 0.72 11.425 1.62 11.405 1.62 11.405 2.01 11.285 2.01 11.285 1.5 10.705 1.5 10.705 1.16 9.765 1.16 9.765 1.04 10.825 1.04 10.825 1.38 11.305 1.38 11.305 0.72 11.225 0.72 11.225 0.6 11.465 0.6 ;
      POLYGON 10.585 1.4 10.04 1.4 10.04 1.77 9.8 1.77 9.8 1.6 9.92 1.6 9.92 1.4 8.205 1.4 8.205 1.77 8.085 1.77 8.085 1.28 8.165 1.28 8.165 0.5 8.285 0.5 8.285 0.74 9.165 0.74 9.165 0.6 9.405 0.6 9.405 0.72 9.285 0.72 9.285 0.86 8.285 0.86 8.285 1.28 10.585 1.28 ;
      POLYGON 9.765 0.68 9.645 0.68 9.645 0.48 8.985 0.48 8.985 0.62 8.745 0.62 8.745 0.5 8.865 0.5 8.865 0.36 9.765 0.36 ;
      POLYGON 7.865 0.72 7.725 0.72 7.725 1.77 7.605 1.77 7.605 0.96 7.245 0.96 7.245 1.17 5.985 1.17 5.985 0.99 5.505 0.99 5.505 0.56 4.685 0.56 4.685 0.52 4.275 0.52 4.275 1.2 4.155 1.2 4.155 0.4 4.805 0.4 4.805 0.44 5.625 0.44 5.625 0.87 6.105 0.87 6.105 1.05 7.125 1.05 7.125 0.84 7.605 0.84 7.605 0.6 7.745 0.6 7.745 0.48 7.865 0.48 ;
      POLYGON 7.485 0.68 7.005 0.68 7.005 0.93 6.225 0.93 6.225 0.75 6.105 0.75 6.105 0.63 6.345 0.63 6.345 0.81 6.885 0.81 6.885 0.56 7.485 0.56 ;
      POLYGON 7.245 1.64 7.125 1.64 7.125 1.57 6.065 1.57 6.065 1.77 5.945 1.77 5.945 1.45 7.125 1.45 7.125 1.4 7.245 1.4 ;
      POLYGON 6.765 0.69 6.525 0.69 6.525 0.51 5.865 0.51 5.865 0.75 5.745 0.75 5.745 0.39 6.645 0.39 6.645 0.57 6.765 0.57 ;
      POLYGON 6.605 2.25 5.465 2.25 5.465 1.675 4.685 1.675 4.685 0.68 4.965 0.68 4.965 0.8 4.805 0.8 4.805 1.555 5.585 1.555 5.585 2.13 6.605 2.13 ;
      POLYGON 5.105 2.25 4.335 2.25 4.335 1.82 4.395 1.82 4.395 1.44 3.615 1.44 3.615 2.21 3.495 2.21 3.495 1.245 2.875 1.245 2.875 1.125 3.495 1.125 3.495 0.64 3.615 0.64 3.615 1.32 4.395 1.32 4.395 0.64 4.515 0.64 4.515 1.94 4.455 1.94 4.455 2.13 5.105 2.13 ;
  END
END DFFSRHQX8

MACRO AOI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X2 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.98 0.99 5.51 1.11 ;
        RECT 4.075 0.94 5.1 0.99 ;
        RECT 4.13 0.87 5.1 0.99 ;
        RECT 4.01 0.99 4.335 1.09 ;
        RECT 4.01 0.99 4.25 1.11 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.53 0.99 3.83 1.11 ;
        RECT 2.915 0.94 3.175 1.11 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.99 1.96 1.11 ;
        RECT 0.595 0.94 1.62 1.03 ;
        RECT 0.735 0.91 1.62 1.03 ;
        RECT 0.56 0.99 0.855 1.11 ;
    END
  END A0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.71 1.11 4.86 1.58 ;
        RECT 4.71 1.11 4.83 1.61 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.15 1.38 1.65 ;
        RECT 1.23 1.15 1.38 1.62 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.23 3.09 1.41 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8288 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.27 1.56 5.39 2.01 ;
        RECT 4.43 1.73 5.39 1.85 ;
        RECT 1.24 0.63 4.73 0.75 ;
        RECT 4.43 1.53 4.55 2.01 ;
        RECT 2.29 1.53 4.55 1.65 ;
        RECT 2.29 0.63 2.41 1.65 ;
        RECT 2.1 1.175 2.41 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.19 -0.18 5.31 0.64 ;
        RECT 3.79 0.39 4.03 0.51 ;
        RECT 3.79 -0.18 3.91 0.51 ;
        RECT 2.21 0.39 2.45 0.51 ;
        RECT 2.21 -0.18 2.33 0.51 ;
        RECT 0.66 -0.18 0.78 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 1.88 2.01 2.12 2.15 ;
        RECT 1.88 2.01 2 2.79 ;
        RECT 1.04 2.01 1.28 2.15 ;
        RECT 1.04 2.01 1.16 2.79 ;
        RECT 0.26 1.56 0.38 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.81 2.25 2.39 2.25 2.39 2.15 2.27 2.15 2.27 2.01 2.51 2.01 2.51 2.13 3.11 2.13 3.11 2.01 3.35 2.01 3.35 2.13 4.01 2.13 4.01 1.77 4.13 1.77 4.13 2.13 4.85 2.13 4.85 1.97 4.97 1.97 4.97 2.13 5.69 2.13 5.69 1.56 5.81 1.56 ;
      POLYGON 3.71 2.01 3.59 2.01 3.59 1.89 2.87 1.89 2.87 2.01 2.75 2.01 2.75 1.89 1.64 1.89 1.64 2.21 1.52 2.21 1.52 1.89 0.8 1.89 0.8 2.21 0.68 2.21 0.68 1.56 0.8 1.56 0.8 1.77 1.52 1.77 1.52 1.56 1.64 1.56 1.64 1.77 3.71 1.77 ;
  END
END AOI222X2

MACRO OR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.835 1.96 1.15 ;
        RECT 1.655 1.03 1.93 1.18 ;
    END
  END A
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1.175 0.525 1.435 ;
        RECT 0.185 1.26 0.405 1.5 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.02 0.845 1.285 ;
        RECT 0.645 1.165 0.82 1.445 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.24 1.295 1.525 ;
        RECT 0.97 1.405 1.295 1.525 ;
        RECT 0.94 1.465 1.09 1.725 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.355 1.175 2.54 1.435 ;
        RECT 2.355 0.66 2.475 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.935 -0.18 2.055 0.71 ;
        RECT 1.035 -0.18 1.155 0.38 ;
        RECT 0.135 -0.18 0.255 0.9 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.935 1.56 2.055 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.235 1.42 1.535 1.42 1.535 1.965 0.475 1.965 0.475 1.7 0.595 1.7 0.595 1.845 1.415 1.845 1.415 0.9 0.555 0.9 0.555 0.66 0.675 0.66 0.675 0.78 1.455 0.78 1.455 0.66 1.575 0.66 1.575 0.9 1.535 0.9 1.535 1.3 2.235 1.3 ;
  END
END OR4X1

MACRO AOI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X4 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.99 3.435 1.11 ;
        RECT 0.595 0.94 0.855 1.11 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.545 0.94 6.665 1.18 ;
        RECT 5.965 0.99 6.665 1.11 ;
        RECT 6.395 0.94 6.665 1.11 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 0.97 5.025 1.09 ;
        RECT 4.365 0.94 4.625 1.09 ;
        RECT 4.285 0.99 4.525 1.11 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.275 1.23 2.795 1.35 ;
        RECT 2.335 1.23 2.595 1.38 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2416 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.805 1.3 6.925 2.01 ;
        RECT 5.965 1.3 6.925 1.42 ;
        RECT 6.545 0.65 6.785 0.77 ;
        RECT 1.555 0.7 6.665 0.82 ;
        RECT 5.965 1.23 6.085 2.01 ;
        RECT 4.025 1.23 6.085 1.35 ;
        RECT 5.705 0.65 5.945 0.82 ;
        RECT 4.865 0.65 5.105 0.82 ;
        RECT 4.025 0.65 4.265 0.82 ;
        RECT 4.025 0.65 4.145 1.35 ;
        RECT 3.785 0.94 4.145 1.09 ;
        RECT 2.715 0.65 2.955 0.82 ;
        RECT 1.435 0.65 1.675 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 7.025 -0.18 7.145 0.64 ;
        RECT 6.125 0.46 6.365 0.58 ;
        RECT 6.125 -0.18 6.245 0.58 ;
        RECT 5.285 0.46 5.525 0.58 ;
        RECT 5.285 -0.18 5.405 0.58 ;
        RECT 4.445 0.46 4.685 0.58 ;
        RECT 4.445 -0.18 4.565 0.58 ;
        RECT 3.605 0.46 3.845 0.58 ;
        RECT 3.605 -0.18 3.725 0.58 ;
        RECT 2.075 0.46 2.315 0.58 ;
        RECT 2.075 -0.18 2.195 0.58 ;
        RECT 0.855 -0.18 0.975 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 3.555 2.07 3.675 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.345 2.25 3.925 2.25 3.925 1.86 3.805 1.86 3.805 1.74 4.045 1.74 4.045 2.13 4.705 2.13 4.705 1.74 4.825 1.74 4.825 2.13 5.545 2.13 5.545 1.47 5.665 1.47 5.665 2.13 6.385 2.13 6.385 1.54 6.505 1.54 6.505 2.13 7.225 2.13 7.225 1.47 7.345 1.47 ;
      POLYGON 5.245 2.01 5.125 2.01 5.125 1.62 4.405 1.62 4.405 2.01 4.285 2.01 4.285 1.62 3.195 1.62 3.195 2.21 3.075 2.21 3.075 1.62 2.355 1.62 2.355 2.21 2.235 2.21 2.235 1.62 1.515 1.62 1.515 2.21 1.395 2.21 1.395 1.62 0.675 1.62 0.675 2.21 0.555 2.21 0.555 1.5 4.285 1.5 4.285 1.47 4.405 1.47 4.405 1.5 5.125 1.5 5.125 1.47 5.245 1.47 ;
  END
END AOI211X4

MACRO BMXIX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.045 2.11 6.365 2.25 ;
        RECT 6.105 2.1 6.365 2.25 ;
        RECT 5.515 2.11 6.365 2.23 ;
        RECT 5.515 0.95 5.635 2.23 ;
        RECT 5.045 0.95 5.635 1.19 ;
    END
  END X2
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.315 0.68 8.435 2.01 ;
        RECT 7.475 1.025 8.435 1.145 ;
        RECT 7.475 0.885 7.76 1.145 ;
        RECT 7.475 0.68 7.595 2.01 ;
    END
  END PPN
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 2.05 1.62 2.17 ;
        RECT 0.99 1.64 1.11 2.17 ;
        RECT 0.725 1.64 1.11 1.76 ;
        RECT 0.56 1.52 0.855 1.64 ;
        RECT 0.595 1.64 1.11 1.67 ;
        RECT 0.56 1.19 0.68 1.64 ;
        RECT 0.52 1.19 0.68 1.43 ;
    END
  END M0
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.74 2.05 3.56 2.17 ;
        RECT 1.74 1.81 1.86 2.17 ;
        RECT 1.23 1.81 1.86 1.93 ;
        RECT 1.23 1.465 1.38 1.93 ;
        RECT 1.23 1.23 1.35 1.93 ;
        RECT 0.8 1.23 1.35 1.35 ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.995 2.25 1.45 ;
        RECT 2.13 0.98 2.25 1.45 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.96 1.3 4.08 1.42 ;
        RECT 3.96 1.17 4.08 1.42 ;
        RECT 2.915 1.23 3.175 1.38 ;
        RECT 2.96 0.36 3.08 1.43 ;
        RECT 2.46 0.36 3.08 0.48 ;
    END
  END M1
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.735 -0.18 8.855 0.73 ;
        RECT 7.895 -0.18 8.015 0.73 ;
        RECT 7.055 -0.18 7.175 0.92 ;
        RECT 3.88 -0.18 4 0.38 ;
        RECT 2.02 -0.18 2.14 0.86 ;
        RECT 0.68 -0.18 0.8 0.83 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.735 1.36 8.855 2.79 ;
        RECT 7.895 1.36 8.015 2.79 ;
        RECT 6.995 2 7.115 2.79 ;
        RECT 3.66 2.29 3.9 2.79 ;
        RECT 2.24 2.29 2.48 2.79 ;
        RECT 0.84 2.29 1.08 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.315 1.84 6.67 1.84 6.67 1.98 5.875 1.98 5.875 1.99 5.755 1.99 5.755 0.83 5.145 0.83 5.145 0.66 5.385 0.66 5.385 0.71 5.875 0.71 5.875 1.86 6.55 1.86 6.55 1.72 7.195 1.72 7.195 1.04 7.315 1.04 ;
      POLYGON 6.755 1.6 6.635 1.6 6.635 0.98 6.235 0.98 6.235 0.86 6.635 0.86 6.635 0.68 6.755 0.68 ;
      POLYGON 6.425 1.74 6.185 1.74 6.185 1.52 5.995 1.52 5.995 0.59 5.565 0.59 5.565 0.48 4.665 0.48 4.665 1.93 3.92 1.93 3.92 1.69 2.675 1.69 2.675 0.8 2.6 0.8 2.6 0.68 2.84 0.68 2.84 0.8 2.795 0.8 2.795 1.57 4.04 1.57 4.04 1.81 4.545 1.81 4.545 0.36 5.685 0.36 5.685 0.47 6.115 0.47 6.115 1.4 6.425 1.4 ;
      POLYGON 5.395 2.17 3.68 2.17 3.68 1.93 1.98 1.93 1.98 1.69 1.5 1.69 1.5 0.77 1.26 0.77 1.26 0.65 1.62 0.65 1.62 1.57 2.1 1.57 2.1 1.81 3.8 1.81 3.8 2.05 5.275 2.05 5.275 1.46 4.805 1.46 4.805 0.84 4.785 0.84 4.785 0.6 4.905 0.6 4.905 0.72 4.925 0.72 4.925 1.34 5.395 1.34 ;
      POLYGON 4.425 0.9 4.32 0.9 4.32 1.57 4.4 1.57 4.4 1.69 4.16 1.69 4.16 1.57 4.2 1.57 4.2 1.05 3.44 1.05 3.44 1.18 3.32 1.18 3.32 0.93 4.2 0.93 4.2 0.78 4.305 0.78 4.305 0.66 4.425 0.66 ;
      POLYGON 1.86 1.43 1.74 1.43 1.74 0.53 1.14 0.53 1.14 0.99 1.36 0.99 1.36 1.11 1.02 1.11 1.02 1.07 0.4 1.07 0.4 1.55 0.44 1.55 0.44 1.79 0.32 1.79 0.32 1.67 0.28 1.67 0.28 0.95 0.26 0.95 0.26 0.59 0.38 0.59 0.38 0.83 0.4 0.83 0.4 0.95 1.02 0.95 1.02 0.41 1.86 0.41 ;
  END
END BMXIX4

MACRO MX4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4XL 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.795 1.04 0.915 1.44 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.32 0.8 1.725 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3 1.16 3.12 1.655 ;
        RECT 2.97 1.16 3.12 1.625 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 1.52 4.335 1.67 ;
        RECT 4.075 1.33 4.245 1.67 ;
        RECT 4.005 1.33 4.245 1.45 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.6 1.225 4.72 1.515 ;
        RECT 4.365 1.225 4.72 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.525 0.97 5.92 1.135 ;
        RECT 5.525 0.94 5.785 1.135 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.105 1.23 6.365 1.38 ;
        RECT 5.46 1.33 6.345 1.43 ;
        RECT 5.58 1.31 6.365 1.38 ;
        RECT 5.58 1.31 5.7 2.17 ;
        RECT 4.105 2.05 5.7 2.17 ;
        RECT 5.46 1.33 5.7 1.45 ;
        RECT 3.765 2.13 4.225 2.25 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.465 0.255 1.705 ;
        RECT 0.135 0.68 0.255 0.92 ;
        RECT 0.07 1.465 0.22 1.725 ;
        RECT 0.095 0.8 0.215 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 5.84 0.46 6.08 0.58 ;
        RECT 5.96 -0.18 6.08 0.58 ;
        RECT 4.54 -0.18 4.66 0.86 ;
        RECT 3.165 0.68 3.405 0.8 ;
        RECT 3.165 -0.18 3.285 0.8 ;
        RECT 0.555 -0.18 0.675 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 6.02 1.71 6.14 2.79 ;
        RECT 4.345 2.29 4.585 2.79 ;
        RECT 2.865 2.02 2.985 2.79 ;
        RECT 0.555 2 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.605 1.71 6.56 1.71 6.56 1.83 6.44 1.83 6.44 1.59 6.485 1.59 6.485 0.86 6.38 0.86 6.38 0.82 5.6 0.82 5.6 0.56 4.98 0.56 4.98 1.31 5.1 1.31 5.1 1.43 4.86 1.43 4.86 1.105 4.22 1.105 4.22 1.12 3.885 1.12 3.885 1.3 3.6 1.3 3.6 1.42 3.48 1.42 3.48 1.18 3.765 1.18 3.765 0.985 4.86 0.985 4.86 0.44 5.28 0.44 5.28 0.36 5.52 0.36 5.52 0.44 5.72 0.44 5.72 0.7 6.38 0.7 6.38 0.62 6.5 0.62 6.5 0.74 6.605 0.74 ;
      POLYGON 5.38 0.8 5.34 0.8 5.34 1.71 5.2 1.71 5.2 1.93 3.985 1.93 3.985 2.01 3.265 2.01 3.265 1.9 2.475 1.9 2.475 1.34 2.535 1.34 2.535 0.66 2.655 0.66 2.655 1.46 2.595 1.46 2.595 1.78 3.385 1.78 3.385 1.89 3.865 1.89 3.865 1.81 5.08 1.81 5.08 1.59 5.22 1.59 5.22 0.8 5.14 0.8 5.14 0.68 5.38 0.68 ;
      POLYGON 4.02 0.865 3.645 0.865 3.645 1.04 3.36 1.04 3.36 1.54 3.625 1.54 3.625 1.65 3.745 1.65 3.745 1.77 3.505 1.77 3.505 1.66 3.24 1.66 3.24 1.04 2.775 1.04 2.775 0.54 1.835 0.54 1.835 0.66 1.695 0.66 1.695 1.58 1.755 1.58 1.755 1.7 1.515 1.7 1.515 1.58 1.575 1.58 1.575 0.54 1.715 0.54 1.715 0.42 2.895 0.42 2.895 0.92 3.525 0.92 3.525 0.745 3.9 0.745 3.9 0.62 4.02 0.62 ;
      POLYGON 2.415 1.22 2.355 1.22 2.355 2.18 1.035 2.18 1.035 0.8 1.095 0.8 1.095 0.68 1.215 0.68 1.215 0.92 1.155 0.92 1.155 2.06 2.235 2.06 2.235 0.98 2.415 0.98 ;
      POLYGON 2.115 1.94 1.275 1.94 1.275 1.34 1.335 1.34 1.335 0.56 0.915 0.56 0.915 0.92 0.575 0.92 0.575 1.2 0.335 1.2 0.335 1.08 0.455 1.08 0.455 0.8 0.795 0.8 0.795 0.44 1.455 0.44 1.455 1.46 1.395 1.46 1.395 1.82 1.995 1.82 1.995 0.66 2.115 0.66 ;
  END
END MX4XL

MACRO TLATX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX2 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.62 0.68 5.74 2.15 ;
        RECT 5.58 1.175 5.74 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.94 0.885 4.28 1.145 ;
        RECT 3.94 0.68 4.06 2.15 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 1.4 3.465 1.67 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.125 0.895 1.355 ;
        RECT 0.595 1.125 0.855 1.38 ;
    END
  END D
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 6.04 1.5 6.16 2.79 ;
        RECT 5.2 1.5 5.32 2.79 ;
        RECT 4.36 1.5 4.48 2.79 ;
        RECT 3.52 1.79 3.64 2.79 ;
        RECT 2.015 2.08 2.255 2.2 ;
        RECT 2.015 2.08 2.135 2.79 ;
        RECT 0.655 1.82 0.775 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 6.04 -0.18 6.16 0.73 ;
        RECT 5.2 -0.18 5.32 0.73 ;
        RECT 4.36 -0.18 4.48 0.73 ;
        RECT 3.46 -0.18 3.58 0.4 ;
        RECT 2.175 -0.18 2.295 0.4 ;
        RECT 0.555 -0.18 0.795 0.34 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.46 1.36 4.9 1.36 4.9 2.15 4.78 2.15 4.78 0.68 4.9 0.68 4.9 1.24 5.46 1.24 ;
      POLYGON 3.82 1.28 2.775 1.28 2.775 1.54 2.735 1.54 2.735 1.72 2.495 1.72 2.495 1.54 1.815 1.54 1.815 1.42 2.655 1.42 2.655 0.68 2.775 0.68 2.775 1.16 3.82 1.16 ;
      POLYGON 3.28 1.97 3.04 1.97 3.04 1.96 1.895 1.96 1.895 2.12 1.015 2.12 1.015 1.62 0.355 1.62 0.355 1.36 0.475 1.36 0.475 1.5 1.015 1.5 1.015 1.36 1.295 1.36 1.295 0.5 1.695 0.5 1.695 0.4 1.935 0.4 1.935 0.5 2.015 0.5 2.015 0.52 2.415 0.52 2.415 0.44 3.165 0.44 3.165 0.92 3.045 0.92 3.045 0.56 2.535 0.56 2.535 0.64 1.895 0.64 1.895 0.62 1.415 0.62 1.415 1.6 1.135 1.6 1.135 2 1.775 2 1.775 1.84 3.16 1.84 3.16 1.85 3.28 1.85 ;
      POLYGON 2.495 1.3 1.655 1.3 1.655 1.88 1.255 1.88 1.255 1.76 1.535 1.76 1.535 0.74 1.775 0.74 1.775 0.86 1.655 0.86 1.655 1.18 2.495 1.18 ;
      POLYGON 1.175 1.24 1.055 1.24 1.055 1.005 0.235 1.005 0.235 1.74 0.355 1.74 0.355 1.98 0.235 1.98 0.235 1.86 0.115 1.86 0.115 0.8 0.135 0.8 0.135 0.68 0.255 0.68 0.255 0.885 1.175 0.885 ;
  END
END TLATX2

MACRO TBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX8 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 0.94 2.435 1.18 ;
        RECT 0.65 0.99 2.435 1.11 ;
        RECT 1.555 0.99 1.795 1.14 ;
        RECT 0.335 1.315 0.8 1.435 ;
        RECT 0.65 0.99 0.8 1.435 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.615 0.36 5.855 0.48 ;
        RECT 3.435 0.49 5.735 0.61 ;
        RECT 5.615 0.36 5.735 0.61 ;
        RECT 4.395 0.365 4.635 0.61 ;
        RECT 3.675 0.365 3.915 0.61 ;
        RECT 2.555 0.44 3.555 0.56 ;
        RECT 1.095 1.34 2.675 1.46 ;
        RECT 2.555 0.44 2.675 1.46 ;
        RECT 1.175 1.23 1.435 1.46 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.215 0.84 9.015 0.96 ;
        RECT 8.895 0.67 9.015 0.96 ;
        RECT 8.755 0.84 8.875 2.21 ;
        RECT 6.74 1.32 8.875 1.44 ;
        RECT 8.055 0.67 8.175 0.96 ;
        RECT 7.915 1.32 8.035 2.21 ;
        RECT 7.215 0.67 7.335 0.96 ;
        RECT 7.075 1.32 7.195 2.21 ;
        RECT 6.74 1.175 6.89 1.44 ;
        RECT 6.235 1.59 6.86 1.71 ;
        RECT 6.74 0.99 6.86 1.71 ;
        RECT 6.375 0.99 6.86 1.11 ;
        RECT 6.375 0.67 6.495 1.11 ;
        RECT 6.235 1.59 6.355 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 9.315 -0.18 9.435 0.72 ;
        RECT 8.475 -0.18 8.595 0.72 ;
        RECT 7.635 -0.18 7.755 0.72 ;
        RECT 6.795 -0.18 6.915 0.72 ;
        RECT 5.895 0.68 6.135 0.8 ;
        RECT 5.975 -0.18 6.095 0.8 ;
        RECT 4.995 -0.18 5.235 0.37 ;
        RECT 4.035 -0.18 4.275 0.37 ;
        RECT 3.075 -0.18 3.315 0.32 ;
        RECT 2.235 -0.18 2.355 0.81 ;
        RECT 0.775 0.51 1.015 0.63 ;
        RECT 0.775 -0.18 0.895 0.63 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 9.175 1.56 9.295 2.79 ;
        RECT 8.335 1.56 8.455 2.79 ;
        RECT 7.495 1.56 7.615 2.79 ;
        RECT 6.655 1.83 6.775 2.79 ;
        RECT 5.815 1.59 5.935 2.79 ;
        RECT 4.415 2.025 4.655 2.145 ;
        RECT 4.415 2.025 4.535 2.79 ;
        RECT 2.715 2.24 2.955 2.79 ;
        RECT 1.875 1.895 1.995 2.79 ;
        RECT 1.035 1.895 1.155 2.79 ;
        RECT 0.135 1.89 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.575 1.47 5.695 1.47 5.695 2.195 4.775 2.195 4.775 1.905 4.27 1.905 4.27 2.195 3.09 2.195 3.09 2.12 2.295 2.12 2.295 1.76 1.575 1.76 1.575 1.94 1.455 1.94 1.455 1.76 0.675 1.76 0.675 1.94 0.555 1.94 0.555 1.76 0.095 1.76 0.095 0.735 0.135 0.735 0.135 0.615 0.255 0.615 0.255 0.735 0.52 0.735 0.52 0.75 1.195 0.75 1.195 0.68 1.775 0.68 1.775 0.8 1.315 0.8 1.315 0.87 0.4 0.87 0.4 0.855 0.215 0.855 0.215 1.64 2.415 1.64 2.415 2 3.21 2 3.21 2.075 4.15 2.075 4.15 1.785 4.895 1.785 4.895 2.075 5.575 2.075 5.575 1.35 6.455 1.35 6.455 1.23 6.575 1.23 ;
      POLYGON 6.215 1.23 6.095 1.23 6.095 1.04 5.375 1.04 5.375 1.955 5.055 1.955 5.055 1.835 5.255 1.835 5.255 1.665 4.015 1.665 4.015 1.955 3.775 1.955 3.775 1.835 3.895 1.835 3.895 1.545 5.255 1.545 5.255 1.04 3.675 1.04 3.675 0.85 3.555 0.85 3.555 0.73 3.795 0.73 3.795 0.92 4.515 0.92 4.515 0.73 4.755 0.73 4.755 0.92 5.475 0.92 5.475 0.73 5.715 0.73 5.715 0.92 6.215 0.92 ;
      POLYGON 5.135 1.28 3.315 1.28 3.315 1.76 3.435 1.76 3.435 1.88 3.195 1.88 3.195 0.8 2.795 0.8 2.795 0.68 3.315 0.68 3.315 1.16 5.135 1.16 ;
  END
END TBUFX8

MACRO NAND2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.33 3.7 1.725 ;
        RECT 3.58 1.24 3.7 1.725 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.26 2.78 1.38 ;
        RECT 2.335 1.23 2.595 1.38 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1072 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.08 1.5 3.2 2.21 ;
        RECT 0.2 1.5 3.2 1.62 ;
        RECT 2.7 0.65 2.94 0.77 ;
        RECT 0.2 0.7 2.82 0.82 ;
        RECT 2.24 1.5 2.36 2.21 ;
        RECT 1.42 0.65 1.66 0.82 ;
        RECT 1.4 1.5 1.52 2.21 ;
        RECT 0.56 1.5 0.68 2.21 ;
        RECT 0.2 1.23 0.565 1.38 ;
        RECT 0.2 0.7 0.32 1.62 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.4 -0.18 3.52 0.64 ;
        RECT 2.06 0.46 2.3 0.58 ;
        RECT 2.06 -0.18 2.18 0.58 ;
        RECT 0.78 0.46 1.02 0.58 ;
        RECT 0.78 -0.18 0.9 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.5 1.845 3.62 2.79 ;
        RECT 2.66 1.74 2.78 2.79 ;
        RECT 1.82 1.74 1.94 2.79 ;
        RECT 0.98 1.74 1.1 2.79 ;
        RECT 0.14 1.74 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.04 2.21 3.92 2.21 3.92 1.68 3.82 1.68 3.82 1.11 0.44 1.11 0.44 0.99 3.82 0.99 3.82 0.59 3.94 0.59 3.94 1.56 4.04 1.56 ;
  END
END NAND2BX4

MACRO SDFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQXL 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 1.32 0.895 1.625 ;
        RECT 0.65 1.41 0.8 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 1.23 5.865 1.35 ;
        RECT 5.235 1.23 5.495 1.38 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.685 1.245 7.185 1.39 ;
        RECT 6.685 1.21 6.945 1.39 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.445 0.95 7.445 1.07 ;
        RECT 6.975 0.94 7.235 1.09 ;
        RECT 6.585 0.94 7.235 1.07 ;
        RECT 6.585 0.93 6.825 1.07 ;
        RECT 6.445 0.95 6.565 1.39 ;
        RECT 6.225 1.47 6.465 1.59 ;
        RECT 6.345 1.27 6.465 1.59 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 1.32 0.315 1.965 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.44 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.145 -0.18 7.265 0.79 ;
        RECT 5.865 -0.18 5.985 0.79 ;
        RECT 3.695 -0.18 3.935 0.34 ;
        RECT 2.015 -0.18 2.255 0.34 ;
        RECT 0.555 -0.18 0.675 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.085 1.95 7.325 2.07 ;
        RECT 7.085 1.95 7.205 2.79 ;
        RECT 5.725 1.95 5.965 2.07 ;
        RECT 5.725 1.95 5.845 2.79 ;
        RECT 3.695 2.08 3.935 2.2 ;
        RECT 3.695 2.08 3.815 2.79 ;
        RECT 2.095 2.08 2.335 2.2 ;
        RECT 2.095 2.08 2.215 2.79 ;
        RECT 0.615 1.845 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.685 2.01 7.565 2.01 7.565 1.63 6.585 1.63 6.585 1.51 7.565 1.51 7.565 0.55 7.685 0.55 ;
      POLYGON 6.625 0.81 6.325 0.81 6.325 1.15 6.105 1.15 6.105 1.71 6.465 1.71 6.465 1.77 6.545 1.77 6.545 2.01 6.425 2.01 6.425 1.89 6.345 1.89 6.345 1.83 4.935 1.83 4.935 1.59 4.995 1.59 4.995 0.74 5.235 0.74 5.235 0.86 5.115 0.86 5.115 1.71 5.985 1.71 5.985 1.03 6.205 1.03 6.205 0.69 6.505 0.69 6.505 0.55 6.625 0.55 ;
      POLYGON 5.625 0.73 5.385 0.73 5.385 0.62 4.875 0.62 4.875 1.46 4.815 1.46 4.815 1.95 5.545 1.95 5.545 2.07 4.695 2.07 4.695 1.22 4.755 1.22 4.755 0.62 3.195 0.62 3.195 1.24 3.075 1.24 3.075 0.5 4.255 0.5 4.255 0.42 4.495 0.42 4.495 0.5 5.505 0.5 5.505 0.61 5.625 0.61 ;
      POLYGON 4.635 0.86 4.515 0.86 4.515 1.38 4.575 1.38 4.575 1.78 4.455 1.78 4.455 1.5 3.735 1.5 3.735 1.38 3.575 1.38 3.575 1.26 3.855 1.26 3.855 1.38 4.395 1.38 4.395 0.74 4.635 0.74 ;
      POLYGON 4.495 2.16 4.255 2.16 4.255 2.02 4.065 2.02 4.065 1.96 3.39 1.96 3.39 2.02 3.175 2.02 3.175 2.16 2.935 2.16 2.935 2.02 2.475 2.02 2.475 1.96 1.155 1.96 1.155 1.965 1.035 1.965 1.035 0.74 1.275 0.74 1.275 0.86 1.155 0.86 1.155 1.84 2.475 1.84 2.475 1.06 2.715 1.06 2.715 1.18 2.595 1.18 2.595 1.9 3.27 1.9 3.27 1.84 4.185 1.84 4.185 1.9 4.375 1.9 4.375 2.04 4.495 2.04 ;
      POLYGON 4.095 1.26 3.975 1.26 3.975 1.14 3.455 1.14 3.455 1.72 3.215 1.72 3.215 1.6 3.335 1.6 3.335 0.86 3.315 0.86 3.315 0.74 3.555 0.74 3.555 0.86 3.455 0.86 3.455 1.02 4.095 1.02 ;
      POLYGON 2.975 1.78 2.855 1.78 2.855 1.48 2.835 1.48 2.835 0.92 2.675 0.92 2.675 0.68 2.305 0.68 2.305 0.58 1.775 0.58 1.775 0.52 1.635 0.52 1.635 0.4 1.895 0.4 1.895 0.46 2.425 0.46 2.425 0.56 2.795 0.56 2.795 0.8 2.955 0.8 2.955 1.36 2.975 1.36 ;
      POLYGON 2.355 1.26 1.735 1.26 1.735 1.6 1.855 1.6 1.855 1.72 1.615 1.72 1.615 0.92 1.535 0.92 1.535 0.8 1.395 0.8 1.395 0.62 0.915 0.62 0.915 1.2 0.395 1.2 0.395 1.08 0.795 1.08 0.795 0.5 1.515 0.5 1.515 0.68 1.655 0.68 1.655 0.8 1.735 0.8 1.735 1.14 2.355 1.14 ;
  END
END SDFFQXL

MACRO AOI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X2 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.815 0.75 4.935 1.17 ;
        RECT 3 0.75 4.935 0.87 ;
        RECT 3 0.75 3.12 1.17 ;
        RECT 2.97 0.885 3.12 1.145 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.39 0.75 2.51 1.17 ;
        RECT 0.475 0.75 2.51 0.87 ;
        RECT 0.475 0.75 0.595 1.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 0.99 2.25 1.11 ;
        RECT 0.94 0.99 1.09 1.435 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.42 0.99 4.615 1.23 ;
        RECT 4.42 0.99 4.57 1.435 ;
        RECT 3.275 0.99 4.615 1.11 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.495 1.23 3.835 1.44 ;
        RECT 3.495 1.23 3.755 1.465 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.23 1.885 1.435 ;
        RECT 1.465 1.23 1.77 1.46 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.8992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.755 1.56 4.875 2.01 ;
        RECT 3.075 1.585 4.875 1.705 ;
        RECT 3.915 1.56 4.035 2.01 ;
        RECT 1.53 0.51 3.995 0.63 ;
        RECT 3.075 1.55 3.195 2.01 ;
        RECT 2.625 1.55 3.195 1.67 ;
        RECT 2.625 1.52 2.885 1.67 ;
        RECT 2.73 0.51 2.85 1.67 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.915 0.46 5.155 0.58 ;
        RECT 4.915 -0.18 5.035 0.58 ;
        RECT 2.65 -0.18 2.89 0.39 ;
        RECT 0.275 0.46 0.515 0.58 ;
        RECT 0.275 -0.18 0.395 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 2.175 2.03 2.415 2.15 ;
        RECT 2.175 2.03 2.295 2.79 ;
        RECT 1.335 2.03 1.575 2.15 ;
        RECT 1.335 2.03 1.455 2.79 ;
        RECT 0.495 2.03 0.735 2.15 ;
        RECT 0.495 2.03 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.295 2.25 2.655 2.25 2.655 1.91 1.935 1.91 1.935 2.21 1.815 2.21 1.815 1.91 1.095 1.91 1.095 2.21 0.975 2.21 0.975 1.91 0.255 1.91 0.255 2.21 0.135 2.21 0.135 1.56 0.255 1.56 0.255 1.79 0.975 1.79 0.975 1.56 1.095 1.56 1.095 1.79 1.815 1.79 1.815 1.58 1.935 1.58 1.935 1.79 2.775 1.79 2.775 2.13 3.495 2.13 3.495 1.825 3.615 1.825 3.615 2.13 4.335 2.13 4.335 1.825 4.455 1.825 4.455 2.13 5.175 2.13 5.175 1.56 5.295 1.56 ;
  END
END AOI33X2

MACRO XNOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2XL 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 0.98 0.87 1.34 ;
        RECT 0.65 1.08 0.8 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.24 2.815 1.36 ;
        RECT 2.045 1.23 2.305 1.38 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.62 0.295 0.885 ;
        RECT 0.135 0.765 0.255 1.76 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.415 0.68 2.655 0.8 ;
        RECT 2.495 -0.18 2.615 0.8 ;
        RECT 0.595 -0.18 0.715 0.86 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.395 2.22 2.635 2.79 ;
        RECT 0.615 2.16 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.055 2 1.995 2 1.995 2.18 1.175 2.18 1.175 2.06 1.875 2.06 1.875 1.88 2.935 1.88 2.935 1.11 1.795 1.11 1.795 1.2 1.675 1.2 1.675 0.96 1.795 0.96 1.795 0.99 2.895 0.99 2.895 0.62 3.015 0.62 3.015 0.87 3.055 0.87 ;
      POLYGON 2.375 0.48 1.195 0.48 1.195 0.62 1.135 0.62 1.135 1.58 1.155 1.58 1.155 1.7 0.915 1.7 0.915 1.58 1.015 1.58 1.015 0.5 1.075 0.5 1.075 0.36 2.375 0.36 ;
      POLYGON 1.555 1.94 0.675 1.94 0.675 1.675 0.41 1.675 0.41 1.2 0.53 1.2 0.53 1.555 0.795 1.555 0.795 1.82 1.435 1.82 1.435 0.62 1.555 0.62 ;
  END
END XNOR2XL

MACRO ADDFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.765 0.83 5.99 0.95 ;
        RECT 2.705 0.78 3.965 0.88 ;
        RECT 3.5 0.83 5.99 0.9 ;
        RECT 2.625 0.76 3.62 0.8 ;
        RECT 2.625 0.65 2.885 0.8 ;
        RECT 2.705 0.65 2.825 0.98 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.45 1.07 6.735 1.29 ;
        RECT 6.615 1.05 6.735 1.29 ;
        RECT 6.45 1.07 6.6 1.435 ;
        RECT 3.55 1.07 6.735 1.19 ;
        RECT 2.065 1.1 3.67 1.22 ;
        RECT 1.465 0.98 2.185 1.1 ;
        RECT 1.345 1.06 1.585 1.18 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.865 1.31 6.33 1.43 ;
        RECT 1.825 1.34 3.985 1.46 ;
        RECT 3.205 1.34 3.465 1.67 ;
        RECT 1.825 1.22 1.945 1.46 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 1.315 0.68 2.205 ;
        RECT 0.1 0.835 0.68 0.955 ;
        RECT 0.56 0.665 0.68 0.955 ;
        RECT 0.07 1.315 0.68 1.435 ;
        RECT 0.07 1.175 0.22 1.435 ;
        RECT 0.1 0.835 0.22 1.435 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.275 0.885 7.47 1.145 ;
        RECT 7.275 0.64 7.395 1.38 ;
        RECT 7.175 1.26 7.295 2.21 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.855 -0.18 6.975 0.69 ;
        RECT 4.545 0.35 4.785 0.47 ;
        RECT 4.545 -0.18 4.665 0.47 ;
        RECT 3.705 -0.18 3.825 0.64 ;
        RECT 1.545 -0.18 1.785 0.34 ;
        RECT 0.14 -0.18 0.26 0.715 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.695 2.03 6.935 2.15 ;
        RECT 6.695 2.03 6.815 2.79 ;
        RECT 4.35 2.27 4.59 2.79 ;
        RECT 3.69 2.21 3.81 2.79 ;
        RECT 1.425 2.06 1.545 2.79 ;
        RECT 0.14 1.555 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.155 1.14 6.975 1.14 6.975 1.91 6.015 1.91 6.015 2.09 5.895 2.09 5.895 1.91 5.67 1.91 5.67 1.99 5.43 1.99 5.43 1.87 5.55 1.87 5.55 1.79 6.855 1.79 6.855 0.93 6.615 0.93 6.615 0.63 5.625 0.63 5.625 0.64 5.505 0.64 5.505 0.4 5.625 0.4 5.625 0.51 6.735 0.51 6.735 0.81 6.975 0.81 6.975 1.02 7.155 1.02 ;
      POLYGON 5.77 1.67 5.31 1.67 5.31 2.15 4.05 2.15 4.05 2.09 3.785 2.09 3.785 2.03 2.65 2.03 2.65 1.96 1.665 1.96 1.665 1.94 0.825 1.94 0.825 1.195 0.34 1.195 0.34 1.075 0.825 1.075 0.825 0.5 2.385 0.5 2.385 0.41 3.125 0.41 3.125 0.46 3.245 0.46 3.245 0.58 3.005 0.58 3.005 0.53 2.505 0.53 2.505 0.92 2.385 0.92 2.385 0.62 0.945 0.62 0.945 1.82 1.785 1.82 1.785 1.84 2.385 1.84 2.385 1.66 2.505 1.66 2.505 1.84 2.77 1.84 2.77 1.91 2.99 1.91 2.99 1.79 3.11 1.79 3.11 1.91 3.905 1.91 3.905 1.97 4.17 1.97 4.17 2.03 5.19 2.03 5.19 1.55 5.77 1.55 ;
      POLYGON 5.205 0.71 4.125 0.71 4.125 0.4 4.245 0.4 4.245 0.59 5.085 0.59 5.085 0.4 5.205 0.4 ;
      POLYGON 5.07 1.91 4.83 1.91 4.83 1.85 4.05 1.85 4.05 1.61 4.17 1.61 4.17 1.73 4.95 1.73 4.95 1.79 5.07 1.79 ;
      RECT 1.065 0.74 2.145 0.86 ;
      POLYGON 2.145 1.72 1.905 1.72 1.905 1.7 1.065 1.7 1.065 1.58 2.025 1.58 2.025 1.6 2.145 1.6 ;
  END
END ADDFX1

MACRO SDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX8 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.345 2.775 2.19 ;
        RECT 2.655 0.665 2.775 0.985 ;
        RECT 2.635 0.865 2.755 1.465 ;
        RECT 0.07 1.025 2.755 1.145 ;
        RECT 1.815 0.665 1.935 2.19 ;
        RECT 0.975 0.665 1.095 2.185 ;
        RECT 0.135 0.665 0.255 2.185 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 1.155 5.205 1.38 ;
        RECT 5.085 0.98 5.205 1.38 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.535 1.2 9.655 1.44 ;
        RECT 9.35 1.2 9.655 1.435 ;
        RECT 9.35 1.175 9.5 1.435 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.21 11.115 1.395 ;
        RECT 10.745 1.21 11.005 1.42 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.275 0.97 11.395 1.21 ;
        RECT 11.035 0.94 11.295 1.09 ;
        RECT 10.275 0.97 11.395 1.09 ;
        RECT 10.015 1 10.395 1.12 ;
        RECT 10.015 1 10.135 1.44 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.075 -0.18 11.195 0.82 ;
        RECT 9.795 -0.18 9.915 0.64 ;
        RECT 7.425 -0.18 7.665 0.37 ;
        RECT 5.325 -0.18 5.565 0.38 ;
        RECT 3.915 -0.18 4.035 0.65 ;
        RECT 3.075 -0.18 3.195 0.65 ;
        RECT 2.235 -0.18 2.355 0.655 ;
        RECT 1.395 -0.18 1.515 0.655 ;
        RECT 0.555 -0.18 0.675 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 10.915 1.78 11.035 2.79 ;
        RECT 9.535 1.85 9.655 2.79 ;
        RECT 7.425 2.07 7.665 2.19 ;
        RECT 7.425 2.07 7.545 2.79 ;
        RECT 5.645 2.1 5.765 2.79 ;
        RECT 3.975 1.54 4.095 2.79 ;
        RECT 3.075 1.445 3.195 2.79 ;
        RECT 2.235 1.445 2.355 2.79 ;
        RECT 1.395 1.445 1.515 2.79 ;
        RECT 0.555 1.445 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.635 1.68 11.555 1.68 11.555 1.8 11.435 1.8 11.435 1.66 10.415 1.66 10.415 1.24 10.535 1.24 10.535 1.54 11.515 1.54 11.515 0.85 11.495 0.85 11.495 0.58 11.615 0.58 11.615 0.73 11.635 0.73 ;
      POLYGON 10.555 0.85 10.155 0.85 10.155 0.88 9.895 0.88 9.895 1.56 10.295 1.56 10.295 2.21 10.175 2.21 10.175 1.68 8.985 1.68 8.985 1.76 8.745 1.76 8.745 1.53 8.865 1.53 8.865 0.72 8.785 0.72 8.785 0.6 9.025 0.6 9.025 0.72 8.985 0.72 8.985 1.56 9.775 1.56 9.775 0.76 10.035 0.76 10.035 0.73 10.435 0.73 10.435 0.59 10.555 0.59 ;
      POLYGON 9.435 0.83 9.315 0.83 9.315 0.48 8.665 0.48 8.665 1.15 8.705 1.15 8.705 1.39 8.665 1.39 8.665 1.41 8.625 1.41 8.625 1.88 9.175 1.88 9.175 2.03 9.295 2.03 9.295 2.15 9.055 2.15 9.055 2 8.505 2 8.505 1.29 8.545 1.29 8.545 0.48 8.065 0.48 8.065 0.88 8.145 0.88 8.145 1.12 7.945 1.12 7.945 0.61 7.185 0.61 7.185 0.48 6.705 0.48 6.705 0.97 6.965 0.97 6.965 1.21 6.845 1.21 6.845 1.09 6.585 1.09 6.585 0.36 7.305 0.36 7.305 0.49 7.945 0.49 7.945 0.36 9.435 0.36 ;
      POLYGON 8.425 0.72 8.385 0.72 8.385 1.99 8.265 1.99 8.265 1.36 7.465 1.36 7.465 1.31 7.325 1.31 7.325 1.19 7.585 1.19 7.585 1.24 8.265 1.24 8.265 0.72 8.185 0.72 8.185 0.6 8.425 0.6 ;
      POLYGON 8.225 2.25 7.985 2.25 7.985 1.95 7.045 1.95 7.045 2.23 5.925 2.23 5.925 0.86 4.825 0.86 4.825 1.5 5.245 1.5 5.245 1.74 5.125 1.74 5.125 1.62 4.705 1.62 4.705 0.6 4.965 0.6 4.965 0.74 6.045 0.74 6.045 2.11 6.585 2.11 6.585 1.33 6.425 1.33 6.425 1.21 6.705 1.21 6.705 2.11 6.925 2.11 6.925 1.83 8.105 1.83 8.105 2.13 8.225 2.13 ;
      POLYGON 7.825 1.12 7.705 1.12 7.705 1.07 7.205 1.07 7.205 1.45 7.125 1.45 7.125 1.71 7.005 1.71 7.005 1.33 7.085 1.33 7.085 0.85 6.825 0.85 6.825 0.6 7.065 0.6 7.065 0.73 7.205 0.73 7.205 0.95 7.705 0.95 7.705 0.88 7.825 0.88 ;
      POLYGON 6.465 1.99 6.345 1.99 6.345 1.57 6.185 1.57 6.185 0.62 5.085 0.62 5.085 0.48 4.275 0.48 4.275 1.18 4.155 1.18 4.155 0.36 5.205 0.36 5.205 0.5 6.305 0.5 6.305 1.45 6.465 1.45 ;
      POLYGON 5.725 1.98 4.515 1.98 4.515 2.19 4.395 2.19 4.395 1.42 3.675 1.42 3.675 2.19 3.555 2.19 3.555 1.54 3.495 1.54 3.495 1.225 2.875 1.225 2.875 1.105 3.495 1.105 3.495 0.6 3.615 0.6 3.615 1.3 4.395 1.3 4.395 0.6 4.515 0.6 4.515 1.86 5.605 1.86 5.605 1.13 5.725 1.13 ;
  END
END SDFFHQX8

MACRO MDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX2 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.465 1.335 1.585 ;
        RECT 1.215 1.345 1.335 1.585 ;
        RECT 0.94 1.465 1.09 1.725 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.485 0.96 6.68 1.2 ;
        RECT 6.45 0.885 6.675 1.145 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.9 1.025 8.06 1.48 ;
        RECT 7.94 1 8.06 1.48 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 1.23 8.685 1.38 ;
        RECT 8.425 1.07 8.545 1.38 ;
        RECT 8.34 0.76 8.46 1.19 ;
        RECT 8.22 1.07 8.545 1.19 ;
        RECT 7.3 0.76 8.46 0.88 ;
        RECT 7.54 0.76 7.78 1.09 ;
        RECT 7.04 1 7.42 1.12 ;
        RECT 7.3 0.76 7.42 1.12 ;
        RECT 7.04 1 7.16 1.44 ;
    END
  END S0
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.68 0.675 2.205 ;
        RECT 0.36 1.175 0.675 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.1 -0.18 8.22 0.64 ;
        RECT 6.82 -0.18 6.94 0.64 ;
        RECT 4.43 0.38 4.67 0.5 ;
        RECT 4.55 -0.18 4.67 0.5 ;
        RECT 2.57 -0.18 2.69 0.68 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 7.94 1.84 8.06 2.79 ;
        RECT 6.56 1.56 6.68 2.79 ;
        RECT 4.43 2.06 4.67 2.18 ;
        RECT 4.43 2.06 4.55 2.79 ;
        RECT 2.31 2.06 2.43 2.79 ;
        RECT 0.975 1.845 1.095 2.79 ;
        RECT 0.135 1.555 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.925 1.72 8.54 1.72 8.54 1.84 8.42 1.84 8.42 1.72 7.44 1.72 7.44 1.24 7.56 1.24 7.56 1.6 8.805 1.6 8.805 0.95 8.58 0.95 8.58 0.59 8.7 0.59 8.7 0.83 8.925 0.83 ;
      POLYGON 7.58 0.64 7.18 0.64 7.18 0.88 6.92 0.88 6.92 1.56 7.32 1.56 7.32 2.21 7.2 2.21 7.2 1.68 6.8 1.68 6.8 1.44 5.99 1.44 5.99 1.58 5.95 1.58 5.95 1.7 5.83 1.7 5.83 1.46 5.87 1.46 5.87 0.72 5.83 0.72 5.83 0.6 6.07 0.6 6.07 0.72 5.99 0.72 5.99 1.32 6.8 1.32 6.8 0.76 7.06 0.76 7.06 0.52 7.46 0.52 7.46 0.4 7.58 0.4 ;
      POLYGON 6.46 0.66 6.34 0.66 6.34 0.48 5.71 0.48 5.71 1.1 5.75 1.1 5.75 1.34 5.71 1.34 5.71 1.91 6.26 1.91 6.26 2.03 5.59 2.03 5.59 0.48 5.11 0.48 5.11 0.92 5.23 0.92 5.23 1.04 4.99 1.04 4.99 0.74 4.19 0.74 4.19 0.48 3.71 0.48 3.71 0.98 3.57 0.98 3.57 1.26 2.99 1.26 2.99 1.38 2.87 1.38 2.87 1.14 3.45 1.14 3.45 0.86 3.59 0.86 3.59 0.36 4.31 0.36 4.31 0.62 4.99 0.62 4.99 0.36 6.46 0.36 ;
      POLYGON 5.47 1.98 5.35 1.98 5.35 1.3 4.29 1.3 4.29 1.18 5.35 1.18 5.35 0.72 5.23 0.72 5.23 0.6 5.47 0.6 ;
      POLYGON 5.25 2.24 5.01 2.24 5.01 1.94 3.89 1.94 3.89 2.22 2.71 2.22 2.71 1.94 2.035 1.94 2.035 1.965 1.515 1.965 1.515 2.085 1.395 2.085 1.395 1.845 1.455 1.845 1.455 0.68 1.575 0.68 1.575 1.845 1.915 1.845 1.915 1.82 2.83 1.82 2.83 2.1 3.77 2.1 3.77 1.22 3.81 1.22 3.81 1.1 3.93 1.1 3.93 1.34 3.89 1.34 3.89 1.82 5.13 1.82 5.13 2.12 5.25 2.12 ;
      POLYGON 4.87 1.06 4.17 1.06 4.17 1.58 4.13 1.58 4.13 1.7 4.01 1.7 4.01 1.46 4.05 1.46 4.05 0.98 3.83 0.98 3.83 0.6 4.07 0.6 4.07 0.86 4.17 0.86 4.17 0.94 4.87 0.94 ;
      POLYGON 3.47 0.72 2.93 0.72 2.93 1.02 2.75 1.02 2.75 1.5 3.11 1.5 3.11 1.46 3.23 1.46 3.23 1.98 3.11 1.98 3.11 1.62 2.07 1.62 2.07 1.34 2.05 1.34 2.05 1.1 2.19 1.1 2.19 1.5 2.63 1.5 2.63 0.9 2.81 0.9 2.81 0.6 3.47 0.6 ;
      POLYGON 2.51 1.38 2.39 1.38 2.39 0.98 1.93 0.98 1.93 1.46 1.95 1.46 1.95 1.7 1.83 1.7 1.83 1.58 1.81 1.58 1.81 0.56 1.335 0.56 1.335 1.18 0.795 1.18 0.795 1.06 1.215 1.06 1.215 0.44 2.27 0.44 2.27 0.86 2.51 0.86 ;
  END
END MDFFHQX2

MACRO DFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX2 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.085 1.1 2.325 1.29 ;
        RECT 2.1 1.1 2.25 1.47 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.725 2.13 7.185 2.25 ;
        RECT 6.725 1.7 6.845 2.25 ;
        RECT 5.925 1.7 6.845 1.82 ;
        RECT 4.305 2.13 6.045 2.25 ;
        RECT 5.925 1.7 6.045 2.25 ;
        RECT 4.305 1.66 4.425 2.25 ;
        RECT 3.52 1.66 4.425 1.78 ;
        RECT 2.725 1.89 3.64 2.01 ;
        RECT 3.52 1.66 3.64 2.01 ;
        RECT 2.625 1.23 2.885 1.38 ;
        RECT 2.725 1.1 2.845 2.01 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 0.94 9.58 1.09 ;
        RECT 9.165 1.08 9.435 1.2 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.51 0.865 10.66 1.32 ;
        RECT 10.51 0.865 10.63 1.34 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.81 0.855 1.96 ;
        RECT 0.555 1.6 0.715 1.96 ;
        RECT 0.555 0.68 0.675 2.21 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.755 -0.18 10.875 0.745 ;
        RECT 9.405 -0.18 9.645 0.34 ;
        RECT 7.805 0.5 8.045 0.62 ;
        RECT 7.805 -0.18 7.925 0.62 ;
        RECT 2.345 0.62 2.585 0.74 ;
        RECT 2.345 -0.18 2.465 0.74 ;
        RECT 0.975 -0.18 1.095 0.82 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.69 1.46 10.81 2.79 ;
        RECT 9.385 1.58 9.505 2.79 ;
        RECT 7.805 2.03 7.925 2.79 ;
        RECT 7.685 2.03 7.925 2.15 ;
        RECT 6.285 1.94 6.405 2.79 ;
        RECT 6.165 1.94 6.405 2.06 ;
        RECT 3.825 1.9 4.065 2.02 ;
        RECT 3.825 1.9 3.945 2.79 ;
        RECT 2.125 1.83 2.365 1.95 ;
        RECT 2.165 1.83 2.285 2.79 ;
        RECT 0.975 1.69 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.455 0.745 10.39 0.745 10.39 1.58 10.27 1.58 10.27 0.58 9.175 0.58 9.175 0.96 9.045 0.96 9.045 1.12 8.925 1.12 8.925 0.84 9.055 0.84 9.055 0.48 8.425 0.48 8.425 1.23 8.545 1.23 8.545 1.35 8.305 1.35 8.305 0.86 7.005 0.86 7.005 1.1 5.565 1.1 5.565 0.98 6.885 0.98 6.885 0.74 8.305 0.74 8.305 0.36 9.285 0.36 9.285 0.46 9.765 0.46 9.765 0.36 10.005 0.36 10.005 0.46 10.455 0.46 ;
      POLYGON 10.125 0.82 10.005 0.82 10.005 1.46 9.925 1.46 9.925 1.82 9.805 1.82 9.805 1.46 9.025 1.46 9.025 2.25 8.045 2.25 8.045 1.91 6.965 1.91 6.965 1.58 5.805 1.58 5.805 2.01 4.545 2.01 4.545 1.22 4.385 1.22 4.385 1.1 4.665 1.1 4.665 1.89 5.025 1.89 5.025 0.82 5.145 0.82 5.145 1.89 5.685 1.89 5.685 1.46 7.085 1.46 7.085 1.79 8.165 1.79 8.165 2.13 8.905 2.13 8.905 1.24 9.025 1.24 9.025 1.34 9.885 1.34 9.885 0.7 10.125 0.7 ;
      POLYGON 8.935 0.72 8.785 0.72 8.785 1.7 8.765 1.7 8.765 2.01 8.645 2.01 8.645 1.59 8.065 1.59 8.065 1.1 7.125 1.1 7.125 0.98 8.185 0.98 8.185 1.47 8.665 1.47 8.665 0.6 8.935 0.6 ;
      POLYGON 7.945 1.34 7.445 1.34 7.445 1.67 7.205 1.67 7.205 1.55 7.325 1.55 7.325 1.34 5.565 1.34 5.565 1.77 5.325 1.77 5.325 0.74 5.265 0.74 5.265 0.5 5.385 0.5 5.385 0.62 5.445 0.62 5.445 0.74 6.465 0.74 6.465 0.6 6.765 0.6 6.765 0.72 6.585 0.72 6.585 0.86 5.445 0.86 5.445 1.22 7.945 1.22 ;
      POLYGON 7.185 0.62 6.945 0.62 6.945 0.48 6.345 0.48 6.345 0.62 6.105 0.62 6.105 0.5 6.225 0.5 6.225 0.36 7.065 0.36 7.065 0.5 7.185 0.5 ;
      POLYGON 4.905 1.77 4.785 1.77 4.785 0.98 4.265 0.98 4.265 1.22 3.005 1.22 3.005 0.98 2.105 0.98 2.105 0.48 1.335 0.48 1.335 1.24 1.215 1.24 1.215 0.36 2.225 0.36 2.225 0.86 3.125 0.86 3.125 1.1 4.145 1.1 4.145 0.86 4.785 0.86 4.785 0.5 4.905 0.5 ;
      POLYGON 4.545 0.68 4.425 0.68 4.425 0.74 4.025 0.74 4.025 0.98 3.305 0.98 3.305 0.74 3.185 0.74 3.185 0.62 3.425 0.62 3.425 0.86 3.905 0.86 3.905 0.62 4.305 0.62 4.305 0.56 4.545 0.56 ;
      POLYGON 4.425 1.54 3.205 1.54 3.205 1.77 2.965 1.77 2.965 1.53 3.085 1.53 3.085 1.42 4.425 1.42 ;
      POLYGON 3.785 0.74 3.665 0.74 3.665 0.5 2.945 0.5 2.945 0.74 2.825 0.74 2.825 0.38 3.785 0.38 ;
      POLYGON 3.705 2.25 2.485 2.25 2.485 1.71 1.705 1.71 1.705 0.72 1.865 0.72 1.865 0.6 1.985 0.6 1.985 0.84 1.825 0.84 1.825 1.59 2.605 1.59 2.605 2.13 3.705 2.13 ;
      POLYGON 2.045 2.25 1.395 2.25 1.395 1.8 1.455 1.8 1.455 1.48 0.815 1.48 0.815 1.22 0.935 1.22 0.935 1.36 1.455 1.36 1.455 0.68 1.575 0.68 1.575 1.92 1.515 1.92 1.515 2.13 2.045 2.13 ;
  END
END DFFSRHQX2

MACRO MX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.605 1.185 1.725 ;
        RECT 1.065 1.31 1.185 1.725 ;
        RECT 0.36 1.465 0.51 1.725 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 1.28 0.885 1.485 ;
        RECT 0.65 1.09 0.8 1.485 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.905 1.24 2.305 1.38 ;
        RECT 2.045 1.23 2.305 1.38 ;
        RECT 1.905 1.24 2.025 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.175 2.83 1.435 ;
        RECT 2.425 1.175 2.83 1.295 ;
        RECT 2.425 0.59 2.545 1.62 ;
        RECT 2.405 1.5 2.525 2.21 ;
        RECT 2.345 0.47 2.465 0.71 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.765 -0.18 2.885 0.65 ;
        RECT 1.925 -0.18 2.045 0.71 ;
        RECT 0.625 -0.18 0.745 0.71 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.825 1.56 2.945 2.79 ;
        RECT 1.985 1.85 2.105 2.79 ;
        RECT 0.705 1.97 0.825 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.305 1.1 2.065 1.1 2.065 0.95 1.785 0.95 1.785 2.01 1.525 2.01 1.525 2.03 1.285 2.03 1.285 1.91 1.405 1.91 1.405 1.89 1.665 1.89 1.665 0.95 1.425 0.95 1.425 0.73 1.265 0.73 1.265 0.47 1.385 0.47 1.385 0.61 1.545 0.61 1.545 0.83 2.305 0.83 ;
      POLYGON 1.545 1.77 1.425 1.77 1.425 1.19 1.065 1.19 1.065 0.97 0.24 0.97 0.24 1.845 0.405 1.845 0.405 2.09 0.285 2.09 0.285 1.965 0.12 1.965 0.12 0.73 0.205 0.73 0.205 0.47 0.325 0.47 0.325 0.85 1.305 0.85 1.305 1.07 1.545 1.07 ;
  END
END MX2X2

MACRO NAND4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.465 ;
        RECT 0.375 1.01 0.495 1.495 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.02 0.835 1.39 ;
        RECT 0.65 1.07 0.8 1.435 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.545 1.03 5.73 1.435 ;
        RECT 5.545 1.015 5.665 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.085 0.95 7.205 1.4 ;
        RECT 7.03 0.775 7.18 1.205 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9392 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.205 0.605 8.325 0.845 ;
        RECT 8.025 0.725 8.325 0.845 ;
        RECT 7.365 0.775 8.145 0.895 ;
        RECT 7.955 1.56 8.075 2.21 ;
        RECT 7.775 1.56 8.075 1.68 ;
        RECT 2.045 1.555 7.895 1.67 ;
        RECT 7.775 0.775 7.895 1.68 ;
        RECT 2.075 1.56 8.075 1.675 ;
        RECT 7.365 0.605 7.485 0.895 ;
        RECT 7.115 1.555 7.235 2.21 ;
        RECT 6.275 1.555 6.395 2.21 ;
        RECT 5.435 1.555 5.555 2.21 ;
        RECT 4.595 1.555 4.715 2.21 ;
        RECT 3.755 1.555 3.875 2.21 ;
        RECT 2.915 1.555 3.035 2.21 ;
        RECT 2.045 1.52 2.305 1.67 ;
        RECT 2.075 1.52 2.195 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 2.715 0.475 2.955 0.595 ;
        RECT 2.835 -0.18 2.955 0.595 ;
        RECT 1.875 0.475 2.115 0.595 ;
        RECT 1.875 -0.18 1.995 0.595 ;
        RECT 0.555 -0.18 0.675 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.375 1.56 8.495 2.79 ;
        RECT 7.535 1.795 7.655 2.79 ;
        RECT 6.695 1.795 6.815 2.79 ;
        RECT 5.855 1.795 5.975 2.79 ;
        RECT 5.015 1.795 5.135 2.79 ;
        RECT 4.175 1.795 4.295 2.79 ;
        RECT 3.335 1.795 3.455 2.79 ;
        RECT 2.495 1.795 2.615 2.79 ;
        RECT 1.655 1.56 1.775 2.79 ;
        RECT 0.555 1.615 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.745 0.655 8.625 0.655 8.625 0.485 7.905 0.485 7.905 0.655 7.785 0.655 7.785 0.485 7.065 0.485 7.065 0.655 6.945 0.655 6.945 0.485 6.225 0.485 6.225 0.655 6.105 0.655 6.105 0.485 5.385 0.485 5.385 0.655 5.265 0.655 5.265 0.365 8.745 0.365 ;
      POLYGON 6.645 0.895 3.795 0.895 3.795 0.885 3.615 0.885 3.615 0.605 3.735 0.605 3.735 0.765 3.915 0.765 3.915 0.775 4.455 0.775 4.455 0.605 4.575 0.605 4.575 0.775 5.685 0.775 5.685 0.605 5.805 0.605 5.805 0.775 6.525 0.775 6.525 0.605 6.645 0.605 ;
      POLYGON 4.995 0.655 4.875 0.655 4.875 0.485 4.155 0.485 4.155 0.655 4.035 0.655 4.035 0.485 3.375 0.485 3.375 0.595 3.27 0.595 3.27 0.835 2.475 0.835 2.475 0.845 2.355 0.845 2.355 0.835 1.635 0.835 1.635 0.845 1.515 0.845 1.515 0.605 1.635 0.605 1.635 0.715 2.355 0.715 2.355 0.605 2.475 0.605 2.475 0.715 3.15 0.715 3.15 0.595 3.135 0.595 3.135 0.475 3.24 0.475 3.24 0.365 4.995 0.365 ;
      POLYGON 3.675 1.125 1.275 1.125 1.275 0.48 0.915 0.48 0.915 0.89 0.24 0.89 0.24 1.585 0.255 1.585 0.255 2.21 0.135 2.21 0.135 1.705 0.12 1.705 0.12 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.77 0.795 0.77 0.795 0.36 1.395 0.36 1.395 1.005 3.675 1.005 ;
      POLYGON 1.975 1.4 1.155 1.4 1.155 1.52 1.095 1.52 1.095 2.21 0.975 2.21 0.975 1.4 1.035 1.4 1.035 0.6 1.155 0.6 1.155 1.28 1.975 1.28 ;
  END
END NAND4BBX4

MACRO BMXIX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX2 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.23 1.335 1.49 ;
        RECT 0.305 1.23 1.335 1.35 ;
        RECT 0.305 1.23 0.565 1.38 ;
        RECT 0.355 1.23 0.475 1.47 ;
    END
  END M0
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.785 2.11 3.435 2.23 ;
        RECT 1 2.03 2.905 2.15 ;
        RECT 1 1.61 1.12 2.15 ;
        RECT 0.735 1.61 1.12 1.73 ;
        RECT 0.595 1.52 0.975 1.67 ;
        RECT 0.735 1.47 0.975 1.73 ;
    END
  END S
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.18 2.305 1.38 ;
        RECT 1.955 1.255 2.195 1.43 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.755 1.25 3.995 1.37 ;
        RECT 2.975 1.31 3.875 1.43 ;
        RECT 3.205 1.23 3.465 1.43 ;
    END
  END M1
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.16 0.885 6.31 1.145 ;
        RECT 6.1 1.025 6.22 1.45 ;
    END
  END X2
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.785 0.67 6.905 1.025 ;
        RECT 6.78 0.885 6.9 1.99 ;
        RECT 6.74 0.885 6.9 1.145 ;
    END
  END PPN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 7.205 -0.18 7.325 0.72 ;
        RECT 6.245 -0.18 6.485 0.37 ;
        RECT 3.555 -0.18 3.795 0.32 ;
        RECT 1.935 -0.18 2.055 0.85 ;
        RECT 0.555 -0.18 0.675 0.85 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 7.2 1.34 7.32 2.79 ;
        RECT 6.36 1.53 6.48 2.79 ;
        RECT 3.555 2.29 3.795 2.79 ;
        RECT 1.995 2.27 2.235 2.79 ;
        RECT 0.715 1.85 0.835 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.62 1.23 6.5 1.23 6.5 0.61 5.705 0.61 5.705 0.51 5.135 0.51 5.135 1.77 5.015 1.77 5.015 0.39 5.825 0.39 5.825 0.49 6.62 0.49 ;
      POLYGON 6.12 1.71 5.795 1.71 5.795 2.25 4.875 2.25 4.875 2.13 5.675 2.13 5.675 1.23 5.495 1.23 5.495 0.99 5.765 0.99 5.765 0.73 6.005 0.73 6.005 0.85 5.885 0.85 5.885 1.11 5.795 1.11 5.795 1.59 6.12 1.59 ;
      POLYGON 5.555 0.87 5.375 0.87 5.375 1.65 5.555 1.65 5.555 2.01 4.755 2.01 4.755 2.17 3.555 2.17 3.555 1.99 3.025 1.99 3.025 1.91 2.695 1.91 2.695 1.79 3.145 1.79 3.145 1.87 3.675 1.87 3.675 2.05 4.635 2.05 4.635 1.89 4.775 1.89 4.775 0.51 4.415 0.51 4.415 0.56 3.3 0.56 3.3 0.61 3.035 0.61 3.035 0.85 2.915 0.85 2.915 0.49 3.18 0.49 3.18 0.44 4.295 0.44 4.295 0.39 4.895 0.39 4.895 1.89 5.435 1.89 5.435 1.77 5.255 1.77 5.255 0.75 5.435 0.75 5.435 0.63 5.555 0.63 ;
      POLYGON 4.655 0.87 4.515 0.87 4.515 1.53 4.655 1.53 4.655 1.77 4.515 1.77 4.515 1.93 3.795 1.93 3.795 1.67 1.575 1.67 1.575 1.91 1.295 1.91 1.295 1.79 1.455 1.79 1.455 0.79 1.135 0.79 1.135 0.67 1.575 0.67 1.575 1.55 3.915 1.55 3.915 1.81 4.395 1.81 4.395 0.75 4.535 0.75 4.535 0.63 4.655 0.63 ;
      POLYGON 4.275 0.8 4.235 0.8 4.235 1.57 4.275 1.57 4.275 1.69 4.035 1.69 4.035 1.57 4.115 1.57 4.115 1.11 2.615 1.11 2.615 1.41 2.495 1.41 2.495 0.99 4.115 0.99 4.115 0.8 4.035 0.8 4.035 0.68 4.275 0.68 ;
      POLYGON 1.815 1.41 1.695 1.41 1.695 0.55 1.015 0.55 1.015 0.99 1.235 0.99 1.235 1.11 0.895 1.11 0.895 1.09 0.185 1.09 0.185 1.73 0.415 1.73 0.415 1.97 0.295 1.97 0.295 1.85 0.065 1.85 0.065 0.73 0.135 0.73 0.135 0.61 0.255 0.61 0.255 0.97 0.895 0.97 0.895 0.43 1.815 0.43 ;
  END
END BMXIX2

MACRO AOI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.045 2.54 1.5 ;
        RECT 2.39 1.025 2.51 1.5 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 0.83 2.015 1.195 ;
        RECT 1.81 0.805 1.96 1.165 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.415 1.06 1.635 1.18 ;
        RECT 0.65 1.06 0.8 1.435 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.805 1.515 0.925 ;
        RECT 1.395 0.635 1.515 0.925 ;
        RECT 0.975 1.555 1.095 2.21 ;
        RECT 0.175 1.555 1.095 1.675 ;
        RECT 0.555 0.635 0.675 0.925 ;
        RECT 0.175 0.805 0.295 1.675 ;
        RECT 0.07 1.175 0.295 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.715 -0.18 2.835 0.875 ;
        RECT 1.815 -0.18 1.935 0.685 ;
        RECT 0.975 -0.18 1.095 0.685 ;
        RECT 0.135 -0.18 0.255 0.685 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 1.615 1.56 1.735 2.79 ;
        RECT 0.335 1.795 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.495 1.74 2.15 1.74 2.15 1.435 1.175 1.435 1.175 1.42 1.055 1.42 1.055 1.3 1.295 1.3 1.295 1.315 2.15 1.315 2.15 0.785 2.295 0.785 2.295 0.635 2.415 0.635 2.415 0.905 2.27 0.905 2.27 1.62 2.495 1.62 ;
  END
END AOI2BB1X2

MACRO TBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX6 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.276 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.315 0.94 2.435 1.18 ;
        RECT 0.65 0.99 2.435 1.11 ;
        RECT 1.555 0.99 1.795 1.14 ;
        RECT 0.335 1.315 0.8 1.435 ;
        RECT 0.65 0.99 0.8 1.435 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.72 0.36 5.96 0.48 ;
        RECT 3.515 0.49 5.84 0.61 ;
        RECT 5.72 0.36 5.84 0.61 ;
        RECT 4.5 0.365 4.74 0.61 ;
        RECT 3.78 0.365 4.02 0.61 ;
        RECT 2.555 0.44 3.635 0.56 ;
        RECT 1.095 1.34 2.675 1.46 ;
        RECT 2.555 0.44 2.675 1.46 ;
        RECT 1.175 1.23 1.435 1.46 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0368 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.32 0.84 8.28 0.96 ;
        RECT 8.16 0.67 8.28 0.96 ;
        RECT 8.14 0.84 8.26 2.21 ;
        RECT 6.74 1.32 8.26 1.44 ;
        RECT 7.32 0.67 7.44 0.96 ;
        RECT 7.3 1.32 7.42 2.21 ;
        RECT 6.74 1.175 6.89 1.44 ;
        RECT 6.46 1.59 6.86 1.71 ;
        RECT 6.74 0.99 6.86 1.71 ;
        RECT 6.48 0.99 6.86 1.11 ;
        RECT 6.48 0.67 6.6 1.11 ;
        RECT 6.46 1.59 6.58 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.58 -0.18 8.7 0.72 ;
        RECT 7.74 -0.18 7.86 0.72 ;
        RECT 6.9 -0.18 7.02 0.72 ;
        RECT 6 0.68 6.24 0.8 ;
        RECT 6.08 -0.18 6.2 0.8 ;
        RECT 5.1 -0.18 5.34 0.37 ;
        RECT 4.14 -0.18 4.38 0.37 ;
        RECT 3.18 -0.18 3.42 0.32 ;
        RECT 2.235 -0.18 2.355 0.81 ;
        RECT 0.775 0.51 1.015 0.63 ;
        RECT 0.775 -0.18 0.895 0.63 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.56 1.56 8.68 2.79 ;
        RECT 7.72 1.56 7.84 2.79 ;
        RECT 6.88 1.83 7 2.79 ;
        RECT 6.04 1.59 6.16 2.79 ;
        RECT 4.64 2.025 4.88 2.145 ;
        RECT 4.64 2.025 4.76 2.79 ;
        RECT 2.715 2.24 2.955 2.79 ;
        RECT 1.875 1.895 1.995 2.79 ;
        RECT 1.035 1.895 1.155 2.79 ;
        RECT 0.135 1.89 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.62 1.47 5.825 1.47 5.825 2.195 5 2.195 5 1.905 4.52 1.905 4.52 2.195 3.62 2.195 3.62 2.12 2.295 2.12 2.295 1.76 1.575 1.76 1.575 1.94 1.455 1.94 1.455 1.76 0.675 1.76 0.675 1.94 0.555 1.94 0.555 1.76 0.095 1.76 0.095 0.735 0.135 0.735 0.135 0.615 0.255 0.615 0.255 0.735 0.52 0.735 0.52 0.75 1.195 0.75 1.195 0.68 1.775 0.68 1.775 0.8 1.315 0.8 1.315 0.87 0.4 0.87 0.4 0.855 0.215 0.855 0.215 1.64 2.415 1.64 2.415 2 3.74 2 3.74 2.075 4.4 2.075 4.4 1.785 5.12 1.785 5.12 2.075 5.705 2.075 5.705 1.35 6.5 1.35 6.5 1.23 6.62 1.23 ;
      POLYGON 6.26 1.23 6.14 1.23 6.14 1.04 5.5 1.04 5.5 1.835 5.52 1.835 5.52 1.955 5.28 1.955 5.28 1.835 5.38 1.835 5.38 1.665 4.28 1.665 4.28 1.955 3.96 1.955 3.96 1.835 4.16 1.835 4.16 1.545 5.38 1.545 5.38 1.04 3.78 1.04 3.78 0.85 3.66 0.85 3.66 0.73 3.9 0.73 3.9 0.92 4.62 0.92 4.62 0.73 4.86 0.73 4.86 0.92 5.58 0.92 5.58 0.73 5.82 0.73 5.82 0.92 6.26 0.92 ;
      POLYGON 5.26 1.28 3.395 1.28 3.395 1.76 3.435 1.76 3.435 1.88 3.195 1.88 3.195 1.76 3.275 1.76 3.275 0.8 2.795 0.8 2.795 0.68 3.395 0.68 3.395 1.16 5.26 1.16 ;
  END
END TBUFX6

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.825 0.82 1.24 ;
        RECT 0.65 0.595 0.8 0.995 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.76 0.51 1.215 ;
        RECT 0.38 0.76 0.5 1.24 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.885 1.175 1.205 ;
        RECT 0.94 0.885 1.09 1.21 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5104 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.36 1.515 2.21 ;
        RECT 1.295 0.645 1.415 1.725 ;
        RECT 1.195 0.525 1.315 0.765 ;
        RECT 1.23 1.36 1.515 1.725 ;
        RECT 0.555 1.36 1.515 1.48 ;
        RECT 0.555 1.36 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.22 -0.18 0.34 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.6 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND3X1

MACRO MX3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X4 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.04 2.35 1.245 ;
        RECT 2.1 1.04 2.25 1.435 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.84 0.76 3.99 1.145 ;
        RECT 3.82 1.025 3.94 1.42 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.16 0.79 4.28 1.32 ;
        RECT 4.13 0.79 4.28 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.28 1.145 5.52 1.345 ;
        RECT 5.29 1.07 5.44 1.46 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.58 5.78 1.7 ;
        RECT 5.66 1.44 5.78 1.7 ;
        RECT 5.58 1.465 5.73 1.725 ;
        RECT 5 1.46 5.12 1.7 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.67 1.28 1.79 2.17 ;
        RECT 1.5 0.56 1.79 0.68 ;
        RECT 1.67 0.44 1.79 0.68 ;
        RECT 0.65 1.28 1.79 1.4 ;
        RECT 0.83 0.77 1.62 0.89 ;
        RECT 1.5 0.56 1.62 0.89 ;
        RECT 0.83 0.6 0.95 2.17 ;
        RECT 0.65 1.175 0.95 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.5 -0.18 5.62 0.64 ;
        RECT 4.22 -0.18 4.34 0.64 ;
        RECT 2.09 -0.18 2.21 0.65 ;
        RECT 1.25 -0.18 1.37 0.65 ;
        RECT 0.41 -0.18 0.53 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.44 1.96 5.68 2.08 ;
        RECT 5.44 1.96 5.56 2.79 ;
        RECT 4.08 1.9 4.2 2.79 ;
        RECT 2.09 1.555 2.21 2.79 ;
        RECT 1.25 1.52 1.37 2.79 ;
        RECT 0.41 1.52 0.53 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.1 1.96 5.86 1.96 5.86 1.84 5.9 1.84 5.9 0.95 5.12 0.95 5.12 1.34 4.76 1.34 4.76 1.54 4.64 1.54 4.64 1.22 5 1.22 5 0.76 5.12 0.76 5.12 0.83 5.9 0.83 5.9 0.52 5.92 0.52 5.92 0.4 6.04 0.4 6.04 0.64 6.02 0.64 6.02 1.84 6.1 1.84 ;
      POLYGON 4.98 0.64 4.88 0.64 4.88 1.1 4.52 1.1 4.52 1.66 4.78 1.66 4.78 1.84 4.9 1.84 4.9 1.96 4.66 1.96 4.66 1.78 3.45 1.78 3.45 2.01 3.21 2.01 3.21 1.58 3.49 1.58 3.49 0.84 3.41 0.84 3.41 0.6 3.53 0.6 3.53 0.72 3.61 0.72 3.61 1.66 4.4 1.66 4.4 0.98 4.76 0.98 4.76 0.52 4.86 0.52 4.86 0.4 4.98 0.4 ;
      POLYGON 3.92 0.64 3.8 0.64 3.8 0.48 3.29 0.48 3.29 0.96 3.37 0.96 3.37 1.2 3.29 1.2 3.29 1.46 3.09 1.46 3.09 2.13 3.6 2.13 3.6 1.96 3.84 1.96 3.84 2.08 3.72 2.08 3.72 2.25 2.97 2.25 2.97 1.4 2.71 1.4 2.71 1.16 2.83 1.16 2.83 1.28 3.17 1.28 3.17 0.36 3.92 0.36 ;
      POLYGON 3.05 0.92 2.59 0.92 2.59 1.52 2.85 1.52 2.85 2.17 2.73 2.17 2.73 1.64 2.47 1.64 2.47 0.92 1.98 0.92 1.98 1.1 1.74 1.1 1.74 0.8 2.93 0.8 2.93 0.6 3.05 0.6 ;
  END
END MX3X4

MACRO NAND4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX1 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.925 0.4 1.165 ;
        RECT 0.06 0.885 0.32 1.145 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.77 1.13 2.91 1.44 ;
        RECT 2.625 1.23 2.91 1.415 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.51 0.99 1.67 1.435 ;
        RECT 1.51 0.965 1.635 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 1.2 1.21 1.39 ;
        RECT 0.885 1.23 1.145 1.445 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5364 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.29 1.555 2.27 1.675 ;
        RECT 2.15 0.485 2.27 1.675 ;
        RECT 2.13 1.465 2.25 2.21 ;
        RECT 0.97 0.485 2.27 0.605 ;
        RECT 2.1 1.465 2.25 1.725 ;
        RECT 1.29 1.555 1.41 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.39 -0.18 2.51 0.66 ;
        RECT 0.14 -0.18 0.26 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.55 1.56 2.67 2.79 ;
        RECT 1.71 1.795 1.83 2.79 ;
        RECT 0.87 1.73 0.99 2.79 ;
        RECT 0.14 1.46 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.15 1.8 3.03 1.8 3.03 1.01 2.65 1.01 2.65 1.11 2.39 1.11 2.39 0.99 2.53 0.99 2.53 0.89 2.95 0.89 2.95 0.61 3.07 0.61 3.07 0.77 3.15 0.77 ;
      POLYGON 2.03 1.11 1.79 1.11 1.79 0.845 0.68 0.845 0.68 1.58 0.56 1.58 0.56 0.525 0.68 0.525 0.68 0.725 1.91 0.725 1.91 0.99 2.03 0.99 ;
  END
END NAND4BBX1

MACRO SEDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRXL 0 0 ;
  SIZE 14.21 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 1.15 6.075 1.38 ;
        RECT 5.865 1.04 5.985 1.45 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.045 0.94 8.165 1.2 ;
        RECT 6.905 0.94 8.165 1.06 ;
        RECT 6.905 0.94 7.025 1.33 ;
        RECT 6.685 1.23 6.945 1.38 ;
        RECT 6.825 1.21 7.025 1.33 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.18 7.525 1.45 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.865 1.37 10.105 1.535 ;
        RECT 9.93 1.37 10.08 1.74 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.085 1.18 13.05 1.3 ;
        RECT 12.485 1.18 12.745 1.38 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.41 1.17 13.695 1.29 ;
        RECT 13.575 1.045 13.695 1.29 ;
        RECT 13.41 1.17 13.56 1.435 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 0.68 0.265 0.94 ;
        RECT 0.135 0.82 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.385 0.62 9.505 1.435 ;
        RECT 9.205 1.51 9.475 1.63 ;
        RECT 9.35 1.175 9.475 1.63 ;
        RECT 9.205 1.51 9.325 1.75 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.21 0.18 ;
        RECT 13.435 -0.18 13.555 0.92 ;
        RECT 11.925 0.46 12.165 0.58 ;
        RECT 11.925 -0.18 12.045 0.58 ;
        RECT 11.435 0.43 11.675 0.55 ;
        RECT 11.435 -0.18 11.555 0.55 ;
        RECT 10.315 0.6 10.555 0.72 ;
        RECT 10.435 -0.18 10.555 0.72 ;
        RECT 8.905 -0.18 9.025 0.815 ;
        RECT 7.085 0.46 7.325 0.58 ;
        RECT 7.085 -0.18 7.205 0.58 ;
        RECT 5.725 -0.18 5.845 0.68 ;
        RECT 3.615 0.61 3.855 0.73 ;
        RECT 3.735 -0.18 3.855 0.73 ;
        RECT 1.915 -0.18 2.035 0.86 ;
        RECT 0.565 -0.18 0.685 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.21 2.79 ;
        RECT 13.495 2.08 13.615 2.79 ;
        RECT 10.075 2.23 10.195 2.79 ;
        RECT 8.665 2.25 8.905 2.79 ;
        RECT 7.085 2.29 7.325 2.79 ;
        RECT 5.635 2.29 5.875 2.79 ;
        RECT 3.735 1.81 3.855 2.79 ;
        RECT 3.615 1.81 3.855 1.93 ;
        RECT 1.855 1.94 1.975 2.79 ;
        RECT 0.555 2.16 0.795 2.28 ;
        RECT 0.555 2.16 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.075 1.92 13.28 1.92 13.28 2.18 12.425 2.18 12.425 2.06 13.16 2.06 13.16 1.8 13.955 1.8 13.955 1.68 13.855 1.68 13.855 0.68 13.975 0.68 13.975 1.56 14.075 1.56 ;
      POLYGON 13.29 1.56 13.135 1.56 13.135 1.68 13.015 1.68 13.015 1.44 13.17 1.44 13.17 1.06 11.415 1.06 11.415 1.15 11.295 1.15 11.295 0.91 11.415 0.91 11.415 0.94 12.955 0.94 12.955 0.74 13.195 0.74 13.195 0.94 13.29 0.94 ;
      POLYGON 12.805 0.58 12.42 0.58 12.42 0.82 11.535 0.82 11.535 0.79 11.175 0.79 11.175 1.27 11.905 1.27 11.905 1.44 12.365 1.44 12.365 1.5 12.805 1.5 12.805 1.74 12.565 1.74 12.565 1.62 12.245 1.62 12.245 1.56 11.905 1.56 11.905 1.8 11.785 1.8 11.785 1.39 11.055 1.39 11.055 0.79 10.915 0.79 10.915 0.96 10.075 0.96 10.075 0.48 9.4 0.48 9.4 0.5 9.265 0.5 9.265 1.055 8.885 1.055 8.885 1.12 8.645 1.12 8.645 1 8.765 1 8.765 0.935 9.145 0.935 9.145 0.38 9.28 0.38 9.28 0.36 10.195 0.36 10.195 0.84 10.795 0.84 10.795 0.54 10.915 0.54 10.915 0.66 11.175 0.66 11.175 0.67 11.655 0.67 11.655 0.7 12.3 0.7 12.3 0.46 12.805 0.46 ;
      POLYGON 12.385 1.86 12.265 1.86 12.265 2.04 11.91 2.04 11.91 2.11 10.995 2.11 10.995 1.99 10.975 1.99 10.975 1.75 11.095 1.75 11.095 1.87 11.115 1.87 11.115 1.99 11.79 1.99 11.79 1.92 12.145 1.92 12.145 1.74 12.385 1.74 ;
      POLYGON 11.515 1.87 11.395 1.87 11.395 1.63 10.675 1.63 10.675 1.87 10.555 1.87 10.555 1.51 11.515 1.51 ;
      POLYGON 10.875 2.25 10.37 2.25 10.37 2.11 9.925 2.11 9.925 2.13 8.335 2.13 8.335 2.17 3.975 2.17 3.975 1.69 3.495 1.69 3.495 2.11 2.375 2.11 2.375 2.25 2.135 2.25 2.135 2.13 2.17 2.13 2.17 1.82 1.495 1.82 1.495 1.87 1.375 1.87 1.375 1.82 1.025 1.82 1.025 1.96 0.785 1.96 0.785 1.84 0.905 1.84 0.905 1.7 1.375 1.7 1.375 0.68 1.675 0.68 1.675 0.8 1.495 0.8 1.495 1.7 2.29 1.7 2.29 1.99 3.375 1.99 3.375 1.57 4.095 1.57 4.095 2.05 8.215 2.05 8.215 2.01 9.805 2.01 9.805 1.99 10.49 1.99 10.49 2.13 10.875 2.13 ;
      POLYGON 10.465 1.25 9.745 1.25 9.745 1.675 9.715 1.675 9.715 1.87 9.595 1.87 9.595 1.555 9.625 1.555 9.625 0.6 9.955 0.6 9.955 0.72 9.745 0.72 9.745 1.13 10.465 1.13 ;
      POLYGON 8.525 0.48 7.875 0.48 7.875 0.82 6.785 0.82 6.785 0.86 6.565 0.86 6.565 1.57 7.645 1.57 7.645 1.25 7.885 1.25 7.885 1.37 7.765 1.37 7.765 1.69 6.445 1.69 6.445 0.74 6.665 0.74 6.665 0.62 6.785 0.62 6.785 0.7 7.755 0.7 7.755 0.36 8.525 0.36 ;
      POLYGON 8.405 1.69 8.005 1.69 8.005 1.93 4.795 1.93 4.795 1.67 4.915 1.67 4.915 0.62 5.035 0.62 5.035 1.81 7.885 1.81 7.885 1.57 8.285 1.57 8.285 0.8 8.145 0.8 8.145 0.68 8.405 0.68 ;
      POLYGON 6.325 1.69 6.085 1.69 6.085 1.57 6.195 1.57 6.195 0.92 5.595 0.92 5.595 1.14 5.475 1.14 5.475 0.8 6.195 0.8 6.195 0.68 6.145 0.68 6.145 0.44 6.265 0.44 6.265 0.56 6.315 0.56 6.315 1.57 6.325 1.57 ;
      POLYGON 5.425 0.68 5.355 0.68 5.355 1.57 5.395 1.57 5.395 1.69 5.155 1.69 5.155 1.57 5.235 1.57 5.235 0.5 4.795 0.5 4.795 1.55 4.675 1.55 4.675 0.5 4.095 0.5 4.095 0.97 3.375 0.97 3.375 0.5 2.535 0.5 2.535 1.22 2.595 1.22 2.595 1.34 2.355 1.34 2.355 1.22 2.415 1.22 2.415 0.38 2.935 0.38 2.935 0.36 3.175 0.36 3.175 0.38 3.495 0.38 3.495 0.85 3.975 0.85 3.975 0.38 4.175 0.38 4.175 0.36 4.415 0.36 4.415 0.38 5.425 0.38 ;
      POLYGON 4.555 0.8 4.495 0.8 4.495 1.87 4.375 1.87 4.375 1.21 3.395 1.21 3.395 1.09 4.375 1.09 4.375 0.8 4.315 0.8 4.315 0.68 4.555 0.68 ;
      POLYGON 4.075 1.45 3.255 1.45 3.255 1.87 3.135 1.87 3.135 0.62 3.255 0.62 3.255 1.33 4.075 1.33 ;
      POLYGON 2.895 0.8 2.835 0.8 2.835 1.87 2.715 1.87 2.715 1.58 1.775 1.58 1.775 1.31 1.895 1.31 1.895 1.46 2.715 1.46 2.715 0.8 2.655 0.8 2.655 0.68 2.895 0.68 ;
      POLYGON 1.105 1.58 0.985 1.58 0.985 1.18 0.375 1.18 0.375 1.06 0.985 1.06 0.985 0.68 1.105 0.68 ;
  END
END SEDFFTRXL

MACRO TLATNTSCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX6 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.82 0.565 1.09 ;
        RECT 0.325 0.76 0.565 1.09 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 0.76 1.09 1.205 ;
        RECT 0.925 0.76 1.045 1.23 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.76 1.385 1.25 ;
        RECT 1.23 0.76 1.385 1.22 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1924 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.445 1.19 8.565 2.21 ;
        RECT 8.445 0.405 8.565 1.04 ;
        RECT 6.74 1.19 8.565 1.31 ;
        RECT 8.265 0.92 8.565 1.04 ;
        RECT 7.605 1.04 8.385 1.31 ;
        RECT 7.605 0.405 7.725 2.21 ;
        RECT 6.74 1.175 6.89 1.435 ;
        RECT 6.765 0.405 6.885 2.21 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 8.025 -0.18 8.145 0.92 ;
        RECT 7.185 -0.18 7.305 0.92 ;
        RECT 6.345 -0.18 6.465 0.83 ;
        RECT 4.945 -0.18 5.185 0.32 ;
        RECT 3.355 -0.18 3.595 0.34 ;
        RECT 1.085 -0.18 1.205 0.64 ;
        RECT 0.245 -0.18 0.365 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 8.025 1.43 8.145 2.79 ;
        RECT 7.185 1.43 7.305 2.79 ;
        RECT 6.345 1.77 6.465 2.79 ;
        RECT 5.505 1.77 5.625 2.79 ;
        RECT 4.665 1.56 4.785 2.79 ;
        RECT 3.195 2.18 3.435 2.3 ;
        RECT 3.195 2.18 3.315 2.79 ;
        RECT 0.965 1.61 1.085 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.605 1.28 6.505 1.28 6.505 1.65 6.045 1.65 6.045 2.21 5.925 2.21 5.925 1.65 5.205 1.65 5.205 2.21 5.085 2.21 5.085 1.53 6.385 1.53 6.385 1.16 5.785 1.16 5.785 0.81 5.705 0.81 5.705 0.57 5.825 0.57 5.825 0.69 5.905 0.69 5.905 1.04 6.605 1.04 ;
      POLYGON 6.265 1.4 6.145 1.4 6.145 1.41 5.025 1.41 5.025 1.18 4.305 1.18 4.305 1.5 4.185 1.5 4.185 1.62 4.305 1.62 4.305 2.01 4.065 2.01 4.065 1.5 3.175 1.5 3.175 1.38 4.185 1.38 4.185 1.06 4.465 1.06 4.465 0.68 4.705 0.68 4.705 0.8 4.585 0.8 4.585 1.06 5.025 1.06 5.025 1.05 5.145 1.05 5.145 1.29 6.025 1.29 6.025 1.28 6.265 1.28 ;
      POLYGON 5.665 1.17 5.545 1.17 5.545 1.05 5.465 1.05 5.465 0.93 4.935 0.93 4.935 0.56 4.215 0.56 4.215 0.8 4.075 0.8 4.075 0.92 4.065 0.92 4.065 1.18 3.055 1.18 3.055 1.62 3.795 1.62 3.795 1.7 3.915 1.7 3.915 1.82 3.675 1.82 3.675 1.74 2.935 1.74 2.935 1.18 2.855 1.18 2.855 1.06 3.945 1.06 3.945 0.8 3.955 0.8 3.955 0.68 4.095 0.68 4.095 0.44 5.055 0.44 5.055 0.81 5.585 0.81 5.585 0.93 5.665 0.93 ;
      POLYGON 4.665 1.42 4.545 1.42 4.545 2.25 3.615 2.25 3.615 2.06 2.555 2.06 2.555 1.82 2.375 1.82 2.375 0.86 2.255 0.86 2.255 0.74 2.495 0.74 2.495 1.7 2.675 1.7 2.675 1.94 3.735 1.94 3.735 2.13 4.425 2.13 4.425 1.3 4.665 1.3 ;
      POLYGON 3.975 0.52 3.835 0.52 3.835 0.58 2.735 0.58 2.735 1.3 2.815 1.3 2.815 1.56 2.695 1.56 2.695 1.42 2.615 1.42 2.615 0.58 2.5 0.58 2.5 0.54 1.625 0.54 1.625 1.55 1.685 1.55 1.685 1.67 1.445 1.67 1.445 1.55 1.505 1.55 1.505 0.4 1.625 0.4 1.625 0.42 2.62 0.42 2.62 0.46 3.715 0.46 3.715 0.4 3.975 0.4 ;
      POLYGON 2.255 1.91 1.205 1.91 1.205 1.49 0.505 1.49 0.505 1.67 0.265 1.67 0.265 1.55 0.385 1.55 0.385 1.37 0.685 1.37 0.685 0.64 0.665 0.64 0.665 0.4 0.785 0.4 0.785 0.52 0.805 0.52 0.805 1.37 1.325 1.37 1.325 1.79 2.015 1.79 2.015 0.92 1.895 0.92 1.895 0.68 2.015 0.68 2.015 0.8 2.135 0.8 2.135 1.64 2.255 1.64 ;
  END
END TLATNTSCAX6

MACRO TBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX12 0 0 ;
  SIZE 12.47 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1584 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.3667 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 0.865 1.335 1.105 ;
        RECT 0.535 0.97 1.335 1.09 ;
        RECT 0.595 0.94 0.855 1.09 ;
        RECT 0.535 0.97 0.655 1.23 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.02 1.18 6.995 1.3 ;
        RECT 6.875 1.06 6.995 1.3 ;
        RECT 4.02 1.02 4.175 1.3 ;
        RECT 3.495 0.9 4.14 1.02 ;
        RECT 3.935 1.02 4.175 1.14 ;
        RECT 3.495 0.36 3.615 1.02 ;
        RECT 2.795 0.36 3.615 0.48 ;
        RECT 2.155 0.76 2.915 0.88 ;
        RECT 2.795 0.36 2.915 0.88 ;
        RECT 2.235 0.76 2.475 1.045 ;
        RECT 2.155 0.365 2.275 0.88 ;
        RECT 1.455 0.365 2.275 0.485 ;
        RECT 0.915 1.225 1.575 1.345 ;
        RECT 1.455 0.365 1.575 1.345 ;
        RECT 1.175 1.225 1.435 1.38 ;
        RECT 0.795 1.21 1.035 1.33 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.795 1.44 11.915 2.21 ;
        RECT 11.775 0.59 11.895 0.83 ;
        RECT 11.615 1.44 11.915 1.56 ;
        RECT 11.595 0.71 11.895 0.83 ;
        RECT 7.755 1.32 11.735 1.44 ;
        RECT 11.595 0.71 11.715 1.44 ;
        RECT 10.095 0.76 11.715 0.88 ;
        RECT 10.955 1.32 11.075 2.21 ;
        RECT 10.935 0.59 11.055 0.88 ;
        RECT 10.115 1.32 10.235 2.21 ;
        RECT 10.095 0.59 10.215 0.88 ;
        RECT 9.275 1.32 9.395 2.21 ;
        RECT 9.255 0.59 9.375 0.83 ;
        RECT 9.075 0.71 9.375 0.83 ;
        RECT 9.075 0.71 9.195 1.44 ;
        RECT 8.415 0.76 9.195 0.88 ;
        RECT 8.435 1.32 8.555 2.21 ;
        RECT 8.415 0.59 8.535 0.88 ;
        RECT 7.755 1.175 8.05 1.44 ;
        RECT 7.595 1.54 7.875 1.66 ;
        RECT 7.755 0.71 7.875 1.66 ;
        RECT 7.575 0.71 7.875 0.83 ;
        RECT 7.595 1.54 7.715 2.21 ;
        RECT 7.575 0.59 7.695 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.47 0.18 ;
        RECT 12.195 -0.18 12.315 0.64 ;
        RECT 11.355 -0.18 11.475 0.64 ;
        RECT 10.515 -0.18 10.635 0.64 ;
        RECT 9.675 -0.18 9.795 0.64 ;
        RECT 8.835 -0.18 8.955 0.64 ;
        RECT 7.995 -0.18 8.115 0.64 ;
        RECT 7.155 -0.18 7.275 0.64 ;
        RECT 6.255 0.46 6.495 0.58 ;
        RECT 6.255 -0.18 6.375 0.58 ;
        RECT 5.415 0.46 5.655 0.58 ;
        RECT 5.415 -0.18 5.535 0.58 ;
        RECT 4.575 0.46 4.815 0.58 ;
        RECT 4.575 -0.18 4.695 0.58 ;
        RECT 3.735 0.52 3.975 0.64 ;
        RECT 3.855 -0.18 3.975 0.64 ;
        RECT 2.395 0.52 2.635 0.64 ;
        RECT 2.515 -0.18 2.635 0.64 ;
        RECT 0.715 -0.18 0.835 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.47 2.79 ;
        RECT 12.215 1.56 12.335 2.79 ;
        RECT 11.375 1.56 11.495 2.79 ;
        RECT 10.535 1.56 10.655 2.79 ;
        RECT 9.695 1.56 9.815 2.79 ;
        RECT 8.855 1.56 8.975 2.79 ;
        RECT 8.015 1.56 8.135 2.79 ;
        RECT 7.175 1.9 7.295 2.79 ;
        RECT 5.655 2.015 5.895 2.135 ;
        RECT 5.655 2.015 5.775 2.79 ;
        RECT 4.235 2.225 4.355 2.79 ;
        RECT 3.355 2.225 3.475 2.79 ;
        RECT 2.515 2.225 2.635 2.79 ;
        RECT 1.575 2.23 1.695 2.79 ;
        RECT 0.555 2.03 0.795 2.15 ;
        RECT 0.555 2.03 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.595 1.42 7.475 1.42 7.475 1.78 6.775 1.78 6.775 2.205 6.04 2.205 6.04 1.895 4.715 1.895 4.715 1.865 3.835 1.865 3.835 1.62 3.055 1.62 3.055 1.64 2.815 1.64 2.815 1.62 2.215 1.62 2.215 1.64 1.975 1.64 1.975 1.62 1.275 1.62 1.275 1.67 1.035 1.67 1.035 1.55 1.155 1.55 1.155 1.5 1.695 1.5 1.695 0.605 1.935 0.605 1.935 0.725 1.815 0.725 1.815 1.5 3.255 1.5 3.255 0.72 3.035 0.72 3.035 0.6 3.375 0.6 3.375 1.5 3.955 1.5 3.955 1.745 4.835 1.745 4.835 1.775 6.16 1.775 6.16 2.085 6.655 2.085 6.655 1.66 7.355 1.66 7.355 1.3 7.595 1.3 ;
      POLYGON 7.415 1.15 7.235 1.15 7.235 1.54 6.535 1.54 6.535 1.965 6.415 1.965 6.415 1.54 5.195 1.54 5.195 1.655 4.955 1.655 4.955 1.535 5.075 1.535 5.075 1.42 7.115 1.42 7.115 0.94 6.735 0.94 6.735 0.82 4.26 0.82 4.26 0.725 4.215 0.725 4.215 0.485 4.335 0.485 4.335 0.605 4.38 0.605 4.38 0.7 5.055 0.7 5.055 0.485 5.175 0.485 5.175 0.7 5.895 0.7 5.895 0.48 6.015 0.48 6.015 0.7 6.69 0.7 6.69 0.6 6.735 0.6 6.735 0.48 6.855 0.48 6.855 0.82 7.415 0.82 ;
      RECT 4.795 0.94 6.435 1.06 ;
      POLYGON 5.035 2.245 4.475 2.245 4.475 2.105 1.56 2.105 1.56 1.91 0.255 1.91 0.255 2.14 0.135 2.14 0.135 1.49 0.295 1.49 0.295 0.65 0.415 0.65 0.415 1.61 0.255 1.61 0.255 1.79 1.68 1.79 1.68 1.985 4.595 1.985 4.595 2.125 5.035 2.125 ;
      POLYGON 3.135 1.285 2.055 1.285 2.055 1.38 1.935 1.38 1.935 1.14 2.055 1.14 2.055 1.165 3.135 1.165 ;
  END
END TBUFX12

MACRO SDFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX4 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.08 0.69 2.44 0.81 ;
        RECT 1.995 1.49 2.235 1.61 ;
        RECT 2.08 0.69 2.2 1.61 ;
        RECT 1.23 0.885 2.2 1.005 ;
        RECT 1.26 0.765 1.54 1.005 ;
        RECT 1.42 0.63 1.54 1.005 ;
        RECT 1.035 1.49 1.38 1.61 ;
        RECT 1.26 0.765 1.38 1.61 ;
        RECT 1.23 0.885 1.38 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.98 0.51 1.435 ;
        RECT 0.39 0.93 0.51 1.435 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.715 1.09 6.835 1.33 ;
        RECT 6.135 1.22 6.735 1.34 ;
        RECT 6.615 1.21 6.835 1.33 ;
        RECT 6.135 0.36 6.255 1.34 ;
        RECT 5.055 0.36 6.255 0.48 ;
        RECT 3.735 0.47 5.175 0.59 ;
        RECT 3.935 0.47 4.055 1.1 ;
        RECT 2.94 0.36 3.855 0.48 ;
        RECT 2.68 0.885 3.06 1.125 ;
        RECT 2.94 0.36 3.06 1.125 ;
        RECT 2.68 0.885 2.83 1.145 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.905 0.97 10.025 1.21 ;
        RECT 9.585 0.97 10.025 1.09 ;
        RECT 9.585 0.94 9.845 1.09 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.09 1.02 11.265 1.44 ;
        RECT 11.145 1 11.265 1.44 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.615 1.23 11.875 1.38 ;
        RECT 11.615 1.07 11.765 1.38 ;
        RECT 11.525 0.76 11.645 1.19 ;
        RECT 10.605 0.76 11.645 0.88 ;
        RECT 10.605 0.76 10.845 1.09 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.285 -0.18 11.405 0.64 ;
        RECT 9.685 0.46 9.925 0.58 ;
        RECT 9.685 -0.18 9.805 0.58 ;
        RECT 6.555 -0.18 6.675 0.68 ;
        RECT 4.395 -0.18 4.635 0.35 ;
        RECT 2.68 -0.18 2.8 0.68 ;
        RECT 1.84 -0.18 1.96 0.68 ;
        RECT 1 -0.18 1.12 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.285 1.8 11.405 2.79 ;
        RECT 9.985 1.85 10.105 2.79 ;
        RECT 9.97 1.69 10.09 1.97 ;
        RECT 7.675 2.21 7.915 2.79 ;
        RECT 6.435 2.21 6.675 2.79 ;
        RECT 4.455 2.23 4.575 2.79 ;
        RECT 3.495 2.23 3.615 2.79 ;
        RECT 2.475 1.97 2.715 2.09 ;
        RECT 2.475 1.97 2.595 2.79 ;
        RECT 1.515 1.97 1.755 2.09 ;
        RECT 1.515 1.97 1.635 2.79 ;
        RECT 0.555 1.97 0.795 2.09 ;
        RECT 0.555 1.97 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.115 1.74 11.705 1.74 11.705 1.68 10.85 1.68 10.85 1.42 10.725 1.42 10.725 1.33 10.225 1.33 10.225 0.94 10.345 0.94 10.345 1.21 10.965 1.21 10.965 1.3 10.97 1.3 10.97 1.56 11.995 1.56 11.995 0.95 11.765 0.95 11.765 0.59 11.885 0.59 11.885 0.83 12.115 0.83 ;
      POLYGON 10.73 2.21 10.61 2.21 10.61 1.68 10.485 1.68 10.485 1.57 9.275 1.57 9.275 1.52 9.155 1.52 9.155 1.4 9.345 1.4 9.345 0.53 8.435 0.53 8.435 0.68 8.315 0.68 8.315 0.41 9.465 0.41 9.465 0.7 10.325 0.7 10.325 0.52 10.565 0.52 10.565 0.64 10.445 0.64 10.445 0.82 9.465 0.82 9.465 1.45 10.605 1.45 10.605 1.56 10.73 1.56 ;
      POLYGON 9.865 2.25 8.075 2.25 8.075 2.09 6.15 2.09 6.15 2.19 5.475 2.19 5.475 2.21 5.235 2.21 5.235 2.19 4.705 2.19 4.705 2.11 3.315 2.11 3.315 1.85 0.135 1.85 0.135 1.675 0.12 1.675 0.12 0.69 0.635 0.69 0.635 0.81 0.24 0.81 0.24 1.555 0.255 1.555 0.255 1.73 3.435 1.73 3.435 1.99 4.825 1.99 4.825 2.07 6.03 2.07 6.03 1.97 8.195 1.97 8.195 2.13 9.865 2.13 ;
      POLYGON 9.645 1.97 9.035 1.97 9.035 2.01 8.315 2.01 8.315 1.85 5.535 1.85 5.535 1.32 5.015 1.32 5.015 1.08 5.135 1.08 5.135 1.2 5.535 1.2 5.535 0.92 5.775 0.92 5.775 1.04 5.655 1.04 5.655 1.73 8.315 1.73 8.315 1.16 7.695 1.16 7.695 1.04 8.435 1.04 8.435 1.89 8.915 1.89 8.915 0.65 9.225 0.65 9.225 0.77 9.035 0.77 9.035 1.85 9.525 1.85 9.525 1.73 9.645 1.73 ;
      POLYGON 8.795 1.77 8.555 1.77 8.555 0.92 6.495 0.92 6.495 1.1 6.375 1.1 6.375 0.8 7.895 0.8 7.895 0.54 8.015 0.54 8.015 0.8 8.675 0.8 8.675 1.4 8.795 1.4 ;
      POLYGON 8.195 1.61 7.195 1.61 7.195 1.49 8.075 1.49 8.075 1.34 8.195 1.34 ;
      POLYGON 7.575 1.29 7.455 1.29 7.455 1.37 7.075 1.37 7.075 1.58 6.015 1.58 6.015 1.61 5.775 1.61 5.775 1.49 5.895 1.49 5.895 0.72 5.775 0.72 5.775 0.6 6.015 0.6 6.015 1.46 6.955 1.46 6.955 1.25 7.335 1.25 7.335 1.17 7.575 1.17 ;
      POLYGON 5.595 0.72 5.415 0.72 5.415 0.83 4.895 0.83 4.895 1.44 5.275 1.44 5.275 1.95 5.155 1.95 5.155 1.56 4.775 1.56 4.775 0.83 4.295 0.83 4.295 1.34 3.595 1.34 3.595 1.09 3.715 1.09 3.715 1.22 4.175 1.22 4.175 0.71 5.295 0.71 5.295 0.6 5.595 0.6 ;
      POLYGON 4.655 1.07 4.535 1.07 4.535 1.58 4.095 1.58 4.095 1.87 3.975 1.87 3.975 1.58 3.195 1.58 3.195 1.61 2.955 1.61 2.955 1.58 2.44 1.58 2.44 1.29 2.32 1.29 2.32 1.17 2.56 1.17 2.56 1.46 3.355 1.46 3.355 0.6 3.615 0.6 3.615 0.72 3.475 0.72 3.475 1.46 4.415 1.46 4.415 0.95 4.655 0.95 ;
  END
END SDFFRHQX4

MACRO NAND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XL 0 0 ;
  SIZE 1.16 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.585 1.175 0.8 1.435 ;
        RECT 0.61 1.055 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.36 1.44 ;
        RECT 0.24 1.04 0.36 1.44 ;
        RECT 0.07 1.175 0.22 1.565 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.48 1.555 1.04 1.675 ;
        RECT 0.92 0.8 1.04 1.675 ;
        RECT 0.65 0.68 0.94 0.855 ;
        RECT 0.68 0.8 1.04 0.92 ;
        RECT 0.65 0.595 0.8 0.855 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.16 0.18 ;
        RECT 0.18 -0.18 0.3 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.16 2.79 ;
        RECT 0.905 2.02 1.025 2.79 ;
        RECT 0.135 2.02 0.255 2.79 ;
    END
  END VDD
END NAND2XL

MACRO DFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX1 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1.09 0.87 1.455 ;
        RECT 0.65 1.09 0.87 1.45 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.195 1.205 5.495 1.42 ;
        RECT 5.235 1.18 5.495 1.42 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.295 0.265 2.21 ;
        RECT 0.07 1.175 0.255 1.435 ;
        RECT 0.135 0.68 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.395 0.45 5.635 0.57 ;
        RECT 5.395 -0.18 5.515 0.57 ;
        RECT 3.795 0.41 4.035 0.53 ;
        RECT 3.915 -0.18 4.035 0.53 ;
        RECT 2.015 -0.18 2.135 0.68 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.395 1.54 5.515 2.79 ;
        RECT 3.795 2.09 4.035 2.21 ;
        RECT 3.795 2.09 3.915 2.79 ;
        RECT 1.715 2.01 1.955 2.13 ;
        RECT 1.715 2.01 1.835 2.79 ;
        RECT 0.565 1.85 0.685 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.055 0.78 6.035 0.78 6.035 1.3 5.995 1.3 5.995 1.71 5.875 1.71 5.875 1.18 5.915 1.18 5.915 0.81 5.015 0.81 5.015 0.48 4.535 0.48 4.535 1.1 4.415 1.1 4.415 0.77 3.555 0.77 3.555 0.48 3.075 0.48 3.075 0.98 3.035 0.98 3.035 1.1 3.015 1.1 3.015 1.16 2.455 1.16 2.455 1.39 2.335 1.39 2.335 1.04 2.895 1.04 2.895 0.86 2.955 0.86 2.955 0.36 3.675 0.36 3.675 0.65 4.415 0.65 4.415 0.36 5.135 0.36 5.135 0.69 5.81 0.69 5.81 0.66 5.935 0.66 5.935 0.54 6.055 0.54 ;
      POLYGON 5.795 1.06 5.015 1.06 5.015 1.97 4.475 1.97 4.475 2.13 4.595 2.13 4.595 2.25 4.355 2.25 4.355 1.97 3.255 1.97 3.255 2.23 2.075 2.23 2.075 1.89 1.4 1.89 1.4 1.98 1.105 1.98 1.105 2.1 0.985 2.1 0.985 1.86 0.995 1.86 0.995 1.29 1.035 1.29 1.035 0.68 1.155 0.68 1.155 1.41 1.115 1.41 1.115 1.86 1.28 1.86 1.28 1.77 2.195 1.77 2.195 2.11 3.135 2.11 3.135 1.25 3.275 1.25 3.275 1.13 3.395 1.13 3.395 1.37 3.255 1.37 3.255 1.85 4.895 1.85 4.895 0.93 5.015 0.93 5.015 0.94 5.795 0.94 ;
      POLYGON 4.895 0.72 4.775 0.72 4.775 1.34 4.675 1.34 4.675 1.73 4.555 1.73 4.555 1.37 3.755 1.37 3.755 1.13 3.875 1.13 3.875 1.25 4.555 1.25 4.555 1.22 4.655 1.22 4.655 0.6 4.895 0.6 ;
      POLYGON 4.195 1.13 4.075 1.13 4.075 1.01 3.635 1.01 3.635 1.61 3.495 1.61 3.495 1.73 3.375 1.73 3.375 1.49 3.515 1.49 3.515 1.01 3.195 1.01 3.195 0.6 3.435 0.6 3.435 0.89 4.195 0.89 ;
      POLYGON 2.835 0.72 2.375 0.72 2.375 0.92 2.215 0.92 2.215 1.51 2.575 1.51 2.575 1.47 2.695 1.47 2.695 1.99 2.575 1.99 2.575 1.63 1.595 1.63 1.595 1.37 1.515 1.37 1.515 1.13 1.715 1.13 1.715 1.51 2.095 1.51 2.095 0.8 2.255 0.8 2.255 0.6 2.835 0.6 ;
      POLYGON 1.975 1.39 1.855 1.39 1.855 1.01 1.395 1.01 1.395 1.53 1.475 1.53 1.475 1.65 1.235 1.65 1.235 1.53 1.275 1.53 1.275 0.56 0.915 0.56 0.915 0.97 0.53 0.97 0.53 1.24 0.41 1.24 0.41 0.85 0.795 0.85 0.795 0.44 1.715 0.44 1.715 0.89 1.975 0.89 ;
  END
END DFFHQX1

MACRO TBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX4 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.04 1.14 1.16 ;
        RECT 0.36 0.885 0.51 1.16 ;
        RECT 0.3 1 0.42 1.24 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.555 0.99 2.835 1.11 ;
        RECT 2.715 0.41 2.835 1.11 ;
        RECT 2.075 0.41 2.835 0.53 ;
        RECT 1.26 0.48 2.195 0.6 ;
        RECT 1.26 1.23 1.725 1.38 ;
        RECT 0.56 1.28 1.585 1.4 ;
        RECT 1.26 0.48 1.38 1.4 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.255 1.315 4.375 2.21 ;
        RECT 3.535 0.76 4.335 0.88 ;
        RECT 4.215 0.59 4.335 0.88 ;
        RECT 3.535 1.315 4.375 1.435 ;
        RECT 3.535 1.175 3.7 1.435 ;
        RECT 3.535 0.71 3.655 1.83 ;
        RECT 3.415 1.71 3.535 2.21 ;
        RECT 3.375 0.71 3.655 0.83 ;
        RECT 3.375 0.59 3.495 0.83 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 4.635 -0.18 4.755 0.64 ;
        RECT 3.795 -0.18 3.915 0.64 ;
        RECT 2.955 -0.18 3.075 0.64 ;
        RECT 1.715 -0.18 1.955 0.36 ;
        RECT 0.78 -0.18 0.9 0.71 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 4.675 1.56 4.795 2.79 ;
        RECT 3.775 1.62 4.015 2.15 ;
        RECT 3.775 1.62 3.895 2.79 ;
        RECT 2.915 1.71 3.035 2.79 ;
        RECT 0.975 2.1 1.215 2.22 ;
        RECT 0.975 2.1 1.095 2.79 ;
        RECT 0.135 1.76 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.415 1.59 2.795 1.59 2.795 1.8 2.53 1.8 2.53 2.25 1.615 2.25 1.615 1.98 0.675 1.98 0.675 2.21 0.555 2.21 0.555 1.64 0.06 1.64 0.06 0.645 0.14 0.645 0.14 0.525 0.26 0.525 0.26 0.765 0.18 0.765 0.18 1.52 0.675 1.52 0.675 1.86 1.735 1.86 1.735 2.13 2.41 2.13 2.41 1.68 2.675 1.68 2.675 1.47 3.295 1.47 3.295 1.22 3.415 1.22 ;
      POLYGON 3.075 1.35 2.435 1.35 2.435 1.56 2.255 1.56 2.255 2.01 2.135 2.01 2.135 1.44 2.315 1.44 2.315 0.65 2.595 0.65 2.595 0.77 2.435 0.77 2.435 1.23 2.955 1.23 2.955 0.91 3.075 0.91 ;
      POLYGON 2.195 1.32 1.965 1.32 1.965 1.74 1.455 1.74 1.455 1.62 1.845 1.62 1.845 0.84 1.5 0.84 1.5 0.72 1.965 0.72 1.965 1.2 2.195 1.2 ;
  END
END TBUFX4

MACRO AOI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2XL 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.192 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.545 1.53 2.785 1.65 ;
        RECT 2.565 0.7 2.685 1.65 ;
        RECT 1.55 0.7 2.685 0.82 ;
        RECT 1.52 0.885 1.67 1.145 ;
        RECT 1.55 0.7 1.67 1.145 ;
    END
  END Y
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.265 0.51 1.73 ;
        RECT 0.36 1.235 0.48 1.73 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 0.85 0.855 1.22 ;
        RECT 0.595 0.905 0.855 1.115 ;
    END
  END A0N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.255 0.97 2.445 1.21 ;
        RECT 2 0.94 2.375 1.09 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.885 1.15 3.175 1.38 ;
        RECT 2.885 1 3.005 1.41 ;
    END
  END B0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.825 -0.18 2.945 0.88 ;
        RECT 1.425 -0.18 1.665 0.34 ;
        RECT 0.555 -0.18 0.675 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 1.765 1.58 1.885 2.79 ;
        RECT 0.595 1.97 0.715 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.205 1.76 3.085 1.76 3.085 1.89 2.305 1.89 2.305 1.64 2.005 1.64 2.005 1.46 1.465 1.46 1.465 1.7 1.345 1.7 1.345 1.34 2.125 1.34 2.125 1.52 2.425 1.52 2.425 1.77 2.965 1.77 2.965 1.64 3.205 1.64 ;
      POLYGON 2.205 0.48 2.085 0.48 2.085 0.58 0.915 0.58 0.915 0.66 0.255 0.66 0.255 0.9 0.24 0.9 0.24 1.85 0.295 1.85 0.295 2.09 0.175 2.09 0.175 1.97 0.12 1.97 0.12 0.78 0.135 0.78 0.135 0.54 0.795 0.54 0.795 0.46 1.965 0.46 1.965 0.36 2.205 0.36 ;
      POLYGON 1.4 1.22 1.28 1.22 1.28 1.1 1.155 1.1 1.155 2.09 1.135 2.09 1.135 2.21 1.015 2.21 1.015 1.97 1.035 1.97 1.035 0.72 1.275 0.72 1.275 0.84 1.155 0.84 1.155 0.98 1.4 0.98 ;
  END
END AOI2BB2XL

MACRO SDFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRXL 0 0 ;
  SIZE 13.05 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.23 2.305 1.5 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.855 2.11 7.635 2.23 ;
        RECT 6.855 1.78 6.975 2.23 ;
        RECT 4.415 1.88 6.975 1.9 ;
        RECT 5.655 1.78 6.975 1.9 ;
        RECT 5.175 1.88 5.775 2 ;
        RECT 3.355 1.78 5.295 1.89 ;
        RECT 3.245 1.77 4.535 1.825 ;
        RECT 3.245 1.705 3.475 1.825 ;
        RECT 3.245 1.465 3.41 1.825 ;
        RECT 3.245 0.94 3.365 1.825 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.215 1.28 10.455 1.4 ;
        RECT 10.165 1.52 10.425 1.67 ;
        RECT 10.215 1.28 10.335 1.67 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.52 11.005 1.67 ;
        RECT 10.755 1.29 10.995 1.67 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 1.47 12.455 1.67 ;
        RECT 11.965 1.47 12.455 1.635 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 0.94 12.455 1.09 ;
        RECT 12.265 0.94 12.385 1.24 ;
        RECT 11.365 1 12.385 1.12 ;
        RECT 11.455 0.96 11.575 1.2 ;
        RECT 11.365 1 11.485 1.77 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 0.68 0.265 1.58 ;
        RECT 0.07 0.885 0.265 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 1.51 1.555 1.75 ;
        RECT 1.375 0.63 1.495 0.87 ;
        RECT 1.23 1.465 1.455 1.725 ;
        RECT 1.335 0.75 1.455 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.05 0.18 ;
        RECT 11.955 -0.18 12.075 0.88 ;
        RECT 10.675 -0.18 10.795 0.88 ;
        RECT 9.685 -0.18 9.925 0.34 ;
        RECT 7.815 -0.18 7.935 0.86 ;
        RECT 3.085 -0.18 3.325 0.32 ;
        RECT 1.795 -0.18 1.915 0.87 ;
        RECT 0.565 -0.18 0.685 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.05 2.79 ;
        RECT 12.245 2.03 12.365 2.79 ;
        RECT 10.675 1.97 10.795 2.79 ;
        RECT 9.865 2.12 9.985 2.79 ;
        RECT 7.755 2.29 7.995 2.79 ;
        RECT 6.135 2.26 6.375 2.79 ;
        RECT 4.455 2.26 4.695 2.79 ;
        RECT 3.135 2.25 3.375 2.79 ;
        RECT 1.855 1.63 1.975 2.79 ;
        RECT 0.565 1.46 0.685 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.845 2.09 12.725 2.09 12.725 1.97 12.575 1.97 12.575 1.91 11.705 1.91 11.705 1.51 11.825 1.51 11.825 1.79 12.575 1.79 12.575 0.82 12.345 0.82 12.345 0.7 12.695 0.7 12.695 1.85 12.845 1.85 ;
      POLYGON 11.625 2.15 11.385 2.15 11.385 2.03 11.125 2.03 11.125 1.12 10.435 1.12 10.435 0.58 8.995 0.58 8.995 0.74 9.085 0.74 9.085 1.3 9.175 1.3 9.175 1.86 9.295 1.86 9.295 1.98 9.055 1.98 9.055 1.42 8.965 1.42 8.965 0.86 8.875 0.86 8.875 0.46 10.555 0.46 10.555 1 11.125 1 11.125 0.76 11.215 0.76 11.215 0.7 11.495 0.7 11.495 0.82 11.335 0.82 11.335 0.88 11.245 0.88 11.245 1.91 11.505 1.91 11.505 2.03 11.625 2.03 ;
      POLYGON 10.435 2.03 10.195 2.03 10.195 2 9.925 2 9.925 1.16 9.535 1.16 9.535 1.04 10.075 1.04 10.075 0.7 10.315 0.7 10.315 0.82 10.195 0.82 10.195 1.16 10.045 1.16 10.045 1.88 10.435 1.88 ;
      POLYGON 9.625 2.22 8.215 2.22 8.215 2.14 7.755 2.14 7.755 1.99 7.095 1.99 7.095 1.65 6.695 1.65 6.695 1.36 6.405 1.36 6.405 1.24 6.815 1.24 6.815 1.53 7.215 1.53 7.215 1.87 7.875 1.87 7.875 2.02 8.335 2.02 8.335 2.1 8.815 2.1 8.815 1.66 8.515 1.66 8.515 1.54 8.635 1.54 8.635 1.12 8.605 1.12 8.605 1 8.845 1 8.845 1.12 8.755 1.12 8.755 1.54 8.935 1.54 8.935 2.1 9.505 2.1 9.505 1.6 9.295 1.6 9.295 0.82 9.205 0.82 9.205 0.7 9.445 0.7 9.445 0.82 9.415 0.82 9.415 1.48 9.625 1.48 ;
      POLYGON 8.695 1.98 8.455 1.98 8.455 1.9 8.275 1.9 8.275 1.16 7.175 1.16 7.175 1.04 8.365 1.04 8.365 0.74 8.455 0.74 8.455 0.62 8.575 0.62 8.575 0.86 8.485 0.86 8.485 1.16 8.395 1.16 8.395 1.78 8.575 1.78 8.575 1.86 8.695 1.86 ;
      POLYGON 8.155 1.41 7.455 1.41 7.455 1.63 7.575 1.63 7.575 1.75 7.335 1.75 7.335 1.41 6.935 1.41 6.935 1.04 6.285 1.04 6.285 1.66 5.885 1.66 5.885 1.54 6.165 1.54 6.165 0.62 6.285 0.62 6.285 0.92 6.935 0.92 6.935 0.8 6.975 0.8 6.975 0.62 7.095 0.62 7.095 0.92 7.055 0.92 7.055 1.29 8.155 1.29 ;
      POLYGON 7.515 0.86 7.395 0.86 7.395 0.62 7.215 0.62 7.215 0.5 6.735 0.5 6.735 0.8 6.495 0.8 6.495 0.68 6.615 0.68 6.615 0.38 7.335 0.38 7.335 0.5 7.515 0.5 ;
      POLYGON 6.735 2.19 6.495 2.19 6.495 2.14 6.015 2.14 6.015 2.24 4.925 2.24 4.925 2.14 4.295 2.14 4.295 2.25 4.175 2.25 4.175 2.14 4.13 2.14 4.13 2.13 3.07 2.13 3.07 2.065 2.275 2.065 2.275 1.63 2.425 1.63 2.425 0.87 2.275 0.87 2.275 0.63 2.395 0.63 2.395 0.75 2.545 0.75 2.545 1.75 2.395 1.75 2.395 1.945 3.19 1.945 3.19 2.01 4.295 2.01 4.295 2.02 5.045 2.02 5.045 2.12 5.895 2.12 5.895 2.02 6.615 2.02 6.615 2.07 6.735 2.07 ;
      POLYGON 6.165 0.48 6.045 0.48 6.045 1.28 5.565 1.28 5.565 1.4 5.445 1.4 5.445 1.16 5.925 1.16 5.925 0.36 6.165 0.36 ;
      POLYGON 5.805 1.04 5.325 1.04 5.325 1.52 5.535 1.52 5.535 1.76 5.415 1.76 5.415 1.64 5.205 1.64 5.205 1.28 3.485 1.28 3.485 0.82 3.025 0.82 3.025 1.22 2.905 1.22 2.905 0.7 3.605 0.7 3.605 1.16 5.205 1.16 5.205 0.92 5.685 0.92 5.685 0.62 5.805 0.62 ;
      POLYGON 5.445 0.8 5.085 0.8 5.085 1.04 4.245 1.04 4.245 0.62 4.365 0.62 4.365 0.92 4.965 0.92 4.965 0.68 5.445 0.68 ;
      POLYGON 5.085 1.66 4.845 1.66 4.845 1.65 3.615 1.65 3.615 1.53 4.965 1.53 4.965 1.54 5.085 1.54 ;
      POLYGON 4.845 0.8 4.605 0.8 4.605 0.5 4.125 0.5 4.125 0.72 3.965 0.72 3.965 0.8 3.725 0.8 3.725 0.68 3.845 0.68 3.845 0.6 4.005 0.6 4.005 0.38 4.725 0.38 4.725 0.68 4.845 0.68 ;
      POLYGON 3.885 0.48 3.725 0.48 3.725 0.56 2.785 0.56 2.785 1.34 2.835 1.34 2.835 1.72 2.715 1.72 2.715 1.46 2.665 1.46 2.665 0.56 2.565 0.56 2.565 0.51 2.155 0.51 2.155 1.11 1.815 1.11 1.815 1.15 1.575 1.15 1.575 0.99 2.035 0.99 2.035 0.39 2.685 0.39 2.685 0.44 3.605 0.44 3.605 0.36 3.885 0.36 ;
      POLYGON 1.105 1.58 0.985 1.58 0.985 1.2 0.385 1.2 0.385 1.08 0.985 1.08 0.985 0.68 1.105 0.68 ;
  END
END SDFFNSRXL

MACRO ADDFHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX1 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.585 0.885 7.76 1.145 ;
        RECT 7.585 0.59 7.705 2.21 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 1.32 0.68 2.21 ;
        RECT 0.56 0.67 0.68 0.96 ;
        RECT 0.1 1.32 0.68 1.44 ;
        RECT 0.1 0.84 0.68 0.96 ;
        RECT 0.1 0.84 0.22 1.44 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.5 1.37 6.62 1.61 ;
        RECT 4.745 1.39 6.62 1.51 ;
        RECT 3.16 1.44 4.865 1.54 ;
        RECT 4.36 1.42 6.62 1.51 ;
        RECT 3.16 1.44 4.6 1.56 ;
        RECT 3.16 1.28 3.4 1.56 ;
        RECT 1.99 1.22 3.28 1.34 ;
        RECT 2.915 1.28 3.4 1.38 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.77 1.11 7.085 1.23 ;
        RECT 6.74 1.13 6.89 1.435 ;
        RECT 6.26 1.13 6.89 1.25 ;
        RECT 3.59 1.18 6.38 1.27 ;
        RECT 4.505 1.15 7.085 1.23 ;
        RECT 3.59 1.18 4.625 1.3 ;
        RECT 3.59 1.02 3.83 1.32 ;
        RECT 3.445 1.02 3.83 1.14 ;
        RECT 1.59 0.98 3.565 1.1 ;
        RECT 1.47 1.06 1.71 1.18 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 0.91 6.14 1.03 ;
        RECT 4.075 0.78 4.195 1.06 ;
        RECT 3.685 0.78 4.195 0.9 ;
        RECT 2.89 0.74 3.805 0.86 ;
        RECT 2.915 0.65 3.175 0.86 ;
    END
  END CI
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.045 2.11 7.285 2.23 ;
        RECT 7.045 2.11 7.165 2.79 ;
        RECT 4.74 2.23 4.86 2.79 ;
        RECT 3.72 2.22 3.96 2.79 ;
        RECT 1.67 1.94 1.91 2.79 ;
        RECT 0.14 1.56 0.26 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.045 0.43 7.285 0.55 ;
        RECT 7.045 -0.18 7.165 0.55 ;
        RECT 4.835 0.43 5.075 0.55 ;
        RECT 4.835 -0.18 4.955 0.55 ;
        RECT 3.995 -0.18 4.115 0.64 ;
        RECT 1.67 -0.18 1.91 0.38 ;
        RECT 0.14 -0.18 0.26 0.72 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.465 1.385 7.325 1.385 7.325 1.99 6.12 1.99 6.12 2.21 6 2.21 6 1.99 5.7 1.99 5.7 2.15 5.58 2.15 5.58 1.87 7.205 1.87 7.205 0.79 5.855 0.79 5.855 0.68 5.735 0.68 5.735 0.56 5.975 0.56 5.975 0.67 6.185 0.67 6.185 0.5 6.305 0.5 6.305 0.67 7.325 0.67 7.325 1.265 7.465 1.265 ;
      POLYGON 5.94 1.75 5.46 1.75 5.46 2.11 4.67 2.11 4.67 2.1 3.2 2.1 3.2 2.2 3.08 2.2 3.08 2.1 2.63 2.1 2.63 2.25 2.03 2.25 2.03 1.82 0.95 1.82 0.95 1.2 0.34 1.2 0.34 1.08 0.95 1.08 0.95 0.5 2.63 0.5 2.63 0.41 3.415 0.41 3.415 0.46 3.535 0.46 3.535 0.58 3.295 0.58 3.295 0.53 2.75 0.53 2.75 0.82 2.63 0.82 2.63 0.62 1.07 0.62 1.07 1.7 2.15 1.7 2.15 2.13 2.51 2.13 2.51 1.98 2.69 1.98 2.69 1.5 2.81 1.5 2.81 1.98 3.08 1.98 3.08 1.68 3.2 1.68 3.2 1.98 4.79 1.98 4.79 1.99 5.34 1.99 5.34 1.63 5.94 1.63 ;
      POLYGON 5.495 0.79 4.475 0.79 4.475 0.68 4.355 0.68 4.355 0.56 4.595 0.56 4.595 0.67 5.375 0.67 5.375 0.5 5.495 0.5 ;
      POLYGON 5.22 1.87 5.1 1.87 5.1 1.86 4.2 1.86 4.2 1.74 5.1 1.74 5.1 1.63 5.22 1.63 ;
      RECT 1.19 0.74 2.39 0.86 ;
      POLYGON 2.39 2.01 2.27 2.01 2.27 1.58 1.25 1.58 1.25 1.34 1.37 1.34 1.37 1.46 2.39 1.46 ;
  END
END ADDFHX1

MACRO SDFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX1 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.165 0.915 1.435 ;
        RECT 0.65 1.15 0.8 1.435 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.305 1.23 2.595 1.39 ;
        RECT 2.145 1.19 2.425 1.32 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.305 0.93 7.425 1.17 ;
        RECT 7.03 0.93 7.425 1.05 ;
        RECT 7.03 0.885 7.18 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 1.21 8.885 1.355 ;
        RECT 8.425 1.21 8.685 1.39 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.045 0.97 9.165 1.21 ;
        RECT 7.785 0.97 9.165 1.09 ;
        RECT 8.715 0.94 8.975 1.09 ;
        RECT 7.785 0.97 7.905 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 2.01 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.845 -0.18 8.965 0.82 ;
        RECT 7.305 -0.18 7.425 0.64 ;
        RECT 4.625 -0.18 4.865 0.39 ;
        RECT 2.285 0.39 2.525 0.51 ;
        RECT 2.285 -0.18 2.405 0.51 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.685 1.75 8.805 2.79 ;
        RECT 7.245 2.22 7.365 2.79 ;
        RECT 5.185 2.28 5.425 2.79 ;
        RECT 4.225 2.01 4.345 2.79 ;
        RECT 4.105 2.01 4.345 2.13 ;
        RECT 2.565 1.75 2.685 2.79 ;
        RECT 2.445 1.75 2.685 1.93 ;
        RECT 1.365 2.01 1.605 2.13 ;
        RECT 1.365 2.01 1.485 2.79 ;
        RECT 0.555 1.555 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.405 1.68 9.325 1.68 9.325 1.8 9.205 1.8 9.205 1.63 8.185 1.63 8.185 1.24 8.305 1.24 8.305 1.51 9.285 1.51 9.285 0.85 9.265 0.85 9.265 0.58 9.385 0.58 9.385 0.73 9.405 0.73 ;
      POLYGON 8.325 0.85 7.665 0.85 7.665 1.56 8.065 1.56 8.065 2.21 7.945 2.21 7.945 1.68 7.665 1.68 7.665 1.98 6.475 1.98 6.475 1.3 6.015 1.3 6.015 0.72 5.965 0.72 5.965 0.6 6.205 0.6 6.205 0.72 6.135 0.72 6.135 1.18 6.595 1.18 6.595 1.86 7.545 1.86 7.545 0.73 8.205 0.73 8.205 0.59 8.325 0.59 ;
      POLYGON 7.105 2.22 5.545 2.22 5.545 2.16 4.465 2.16 4.465 1.89 3.505 1.89 3.505 2.23 2.905 2.23 2.905 1.63 2.325 1.63 2.325 1.89 0.975 1.89 0.975 1.555 1.035 1.555 1.035 0.68 1.155 0.68 1.155 1.77 2.205 1.77 2.205 1.51 2.905 1.51 2.905 0.87 3.025 0.87 3.025 2.11 3.385 2.11 3.385 1.27 3.485 1.27 3.485 1.15 3.605 1.15 3.605 1.39 3.505 1.39 3.505 1.77 4.585 1.77 4.585 2.04 5.665 2.04 5.665 2.1 7.105 2.1 ;
      POLYGON 7.045 1.74 6.79 1.74 6.79 1.06 6.255 1.06 6.255 0.94 6.375 0.94 6.375 0.48 5.425 0.48 5.425 0.86 5.585 0.86 5.585 1.1 5.305 1.1 5.305 0.63 4.385 0.63 4.385 0.48 3.905 0.48 3.905 0.92 4.025 0.92 4.025 1.04 3.785 1.04 3.785 0.36 4.505 0.36 4.505 0.51 5.305 0.51 5.305 0.36 6.495 0.36 6.495 0.94 6.79 0.94 6.79 0.59 6.91 0.59 6.91 1.62 7.045 1.62 ;
      POLYGON 6.175 1.94 6.055 1.94 6.055 1.54 5.825 1.54 5.825 1.56 4.505 1.56 4.505 1.11 4.385 1.11 4.385 0.99 4.625 0.99 4.625 1.44 5.705 1.44 5.705 0.72 5.545 0.72 5.545 0.6 5.825 0.6 5.825 1.42 6.175 1.42 ;
      POLYGON 5.755 1.92 4.705 1.92 4.705 1.68 4.945 1.68 4.945 1.8 5.635 1.8 5.635 1.68 5.755 1.68 ;
      POLYGON 5.145 1.32 5.025 1.32 5.025 0.87 4.265 0.87 4.265 1.65 3.625 1.65 3.625 1.53 4.145 1.53 4.145 0.72 4.025 0.72 4.025 0.6 4.265 0.6 4.265 0.75 5.145 0.75 ;
      POLYGON 3.265 1.99 3.145 1.99 3.145 0.75 1.785 0.75 1.785 1.12 1.665 1.12 1.665 0.63 3.145 0.63 3.145 0.54 3.265 0.54 ;
      POLYGON 2.665 1.11 2.545 1.11 2.545 1.07 2.025 1.07 2.025 1.53 2.085 1.53 2.085 1.65 1.845 1.65 1.845 1.53 1.905 1.53 1.905 1.36 1.425 1.36 1.425 0.56 0.915 0.56 0.915 1.03 0.515 1.03 0.515 1.26 0.395 1.26 0.395 0.91 0.795 0.91 0.795 0.44 1.545 0.44 1.545 1.24 1.905 1.24 1.905 0.95 2.545 0.95 2.545 0.87 2.665 0.87 ;
  END
END SDFFRHQX1

MACRO CLKMX2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X3 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.3 1.505 1.42 ;
        RECT 0.465 1.52 1.385 1.64 ;
        RECT 1.265 1.3 1.385 1.64 ;
        RECT 0.465 1.315 0.585 1.64 ;
        RECT 0.36 1.195 0.565 1.435 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.21 1.145 1.4 ;
        RECT 0.705 1.21 1.145 1.365 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.145 1.23 2.595 1.38 ;
        RECT 2.145 1.2 2.265 1.44 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.485 1.315 3.605 2.21 ;
        RECT 2.825 0.77 3.605 0.89 ;
        RECT 3.485 0.59 3.605 0.89 ;
        RECT 2.825 1.315 3.605 1.435 ;
        RECT 2.825 1.175 3.12 1.435 ;
        RECT 2.645 1.5 2.945 1.62 ;
        RECT 2.825 0.65 2.945 1.62 ;
        RECT 2.585 0.65 2.945 0.77 ;
        RECT 2.645 1.5 2.765 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.065 -0.18 3.185 0.64 ;
        RECT 2.225 -0.18 2.345 0.64 ;
        RECT 0.605 -0.18 0.725 0.815 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.065 1.56 3.185 2.79 ;
        RECT 2.225 1.56 2.345 2.79 ;
        RECT 0.765 1.76 1.005 2.15 ;
        RECT 0.765 1.76 0.885 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.685 1.09 2.445 1.09 2.445 1.08 2.025 1.08 2.025 1.68 1.705 1.68 1.705 2.21 1.585 2.21 1.585 1.56 1.905 1.56 1.905 1.08 1.865 1.08 1.865 0.77 1.185 0.77 1.185 0.65 1.985 0.65 1.985 0.96 2.685 0.96 ;
      POLYGON 1.785 1.44 1.665 1.44 1.665 1.32 1.625 1.32 1.625 1.09 1.045 1.09 1.045 1.055 0.24 1.055 0.24 1.555 0.345 1.555 0.345 1.8 0.225 1.8 0.225 1.675 0.12 1.675 0.12 0.815 0.185 0.815 0.185 0.575 0.305 0.575 0.305 0.935 1.745 0.935 1.745 1.2 1.785 1.2 ;
  END
END CLKMX2X3

MACRO EDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX1 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.945 1.1 2.08 1.34 ;
        RECT 1.81 1.175 1.975 1.435 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.56 1.35 7.8 1.52 ;
        RECT 7.61 1.35 7.76 1.725 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.52 10.715 1.67 ;
        RECT 10.455 1.32 10.675 1.67 ;
        RECT 9.795 1.32 10.675 1.44 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.33 1.175 11.53 1.45 ;
        RECT 11.345 1.04 11.515 1.45 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2888 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.38 0.68 1.5 1.025 ;
        RECT 1.33 0.885 1.45 2.21 ;
        RECT 1.23 0.885 1.45 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.255 -0.18 11.375 0.92 ;
        RECT 9.535 0.6 9.775 0.72 ;
        RECT 9.535 -0.18 9.655 0.72 ;
        RECT 8.94 0.6 9.18 0.72 ;
        RECT 8.94 -0.18 9.06 0.72 ;
        RECT 7.88 0.6 8.12 0.72 ;
        RECT 8 -0.18 8.12 0.72 ;
        RECT 6.41 -0.18 6.65 0.32 ;
        RECT 4.81 0.57 5.05 0.69 ;
        RECT 4.81 -0.18 4.93 0.69 ;
        RECT 3.09 0.68 3.33 0.8 ;
        RECT 3.21 -0.18 3.33 0.8 ;
        RECT 1.8 -0.18 1.92 0.92 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.315 1.96 11.435 2.79 ;
        RECT 7.785 2.22 7.905 2.79 ;
        RECT 6.31 2.17 6.55 2.29 ;
        RECT 6.31 2.17 6.43 2.79 ;
        RECT 4.71 2.23 4.83 2.79 ;
        RECT 3.01 1.87 3.27 1.99 ;
        RECT 3.15 1.64 3.27 1.99 ;
        RECT 3.01 1.87 3.13 2.79 ;
        RECT 1.75 2.1 1.99 2.22 ;
        RECT 1.75 2.1 1.87 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.915 1.84 11.12 1.84 11.12 2.15 10.375 2.15 10.375 2.24 10.135 2.24 10.135 2.12 10.255 2.12 10.255 2.03 11 2.03 11 1.72 11.795 1.72 11.795 0.92 11.675 0.92 11.675 0.68 11.795 0.68 11.795 0.8 11.915 0.8 ;
      POLYGON 10.955 1.6 10.835 1.6 10.835 1.2 8.885 1.2 8.885 1.08 10.835 1.08 10.835 0.68 10.955 0.68 ;
      POLYGON 10.515 1.91 10.215 1.91 10.215 1.68 9.615 1.68 9.615 1.86 9.495 1.86 9.495 1.44 8.645 1.44 8.645 0.96 7.64 0.96 7.64 0.48 6.89 0.48 6.89 0.56 6.17 0.56 6.17 0.48 6.05 0.48 6.05 0.36 6.29 0.36 6.29 0.44 6.77 0.44 6.77 0.36 7.76 0.36 7.76 0.84 8.36 0.84 8.36 0.54 8.48 0.54 8.48 0.66 8.765 0.66 8.765 0.84 9.91 0.84 9.91 0.6 10.415 0.6 10.415 0.72 10.03 0.72 10.03 0.96 8.765 0.96 8.765 1.32 9.615 1.32 9.615 1.56 10.335 1.56 10.335 1.79 10.515 1.79 ;
      POLYGON 10.095 1.92 9.975 1.92 9.975 2.1 8.745 2.1 8.745 1.92 8.625 1.92 8.625 1.8 8.865 1.8 8.865 1.98 9.855 1.98 9.855 1.8 10.095 1.8 ;
      POLYGON 9.225 1.86 9.105 1.86 9.105 1.68 8.385 1.68 8.385 1.86 8.265 1.86 8.265 1.56 9.225 1.56 ;
      POLYGON 8.585 2.24 8.345 2.24 8.345 2.1 7.02 2.1 7.02 2.05 6.19 2.05 6.19 2.11 3.51 2.11 3.51 2.25 3.25 2.25 3.25 2.13 3.39 2.13 3.39 1.52 2.85 1.52 2.85 1.99 2.73 1.99 2.73 1.98 1.57 1.98 1.57 1.24 1.69 1.24 1.69 1.86 2.63 1.86 2.63 1.59 2.61 1.59 2.61 0.68 2.73 0.68 2.73 1.4 3.51 1.4 3.51 1.99 6.07 1.99 6.07 1.93 7.14 1.93 7.14 1.98 8.465 1.98 8.465 2.12 8.585 2.12 ;
      POLYGON 8.165 1.23 7.44 1.23 7.44 1.74 7.425 1.74 7.425 1.86 7.305 1.86 7.305 1.62 7.32 1.62 7.32 0.72 7.28 0.72 7.28 0.6 7.52 0.6 7.52 0.72 7.44 0.72 7.44 1.11 8.165 1.11 ;
      POLYGON 7.13 0.8 7.01 0.8 7.01 1.69 7.03 1.69 7.03 1.81 6.79 1.81 6.79 1.69 6.89 1.69 6.89 1.44 5.75 1.44 5.75 1.32 6.89 1.32 6.89 0.68 7.13 0.68 ;
      POLYGON 6.75 1.12 5.79 1.12 5.79 1 5.81 1 5.81 0.5 5.39 0.5 5.39 1.55 5.27 1.55 5.27 0.93 4.57 0.93 4.57 0.5 4.21 0.5 4.21 1.37 4.27 1.37 4.27 1.49 4.03 1.49 4.03 1.37 4.09 1.37 4.09 0.5 3.57 0.5 3.57 1.04 2.85 1.04 2.85 0.56 2.34 0.56 2.34 0.8 2.35 0.8 2.35 1.62 2.47 1.62 2.47 1.74 2.23 1.74 2.23 0.92 2.22 0.92 2.22 0.44 2.97 0.44 2.97 0.92 3.45 0.92 3.45 0.38 3.59 0.38 3.59 0.36 3.83 0.36 3.83 0.38 4.69 0.38 4.69 0.81 5.27 0.81 5.27 0.38 5.93 0.38 5.93 1 6.75 1 ;
      POLYGON 5.69 0.86 5.63 0.86 5.63 1.87 5.51 1.87 5.51 1.79 5.03 1.79 5.03 1.49 4.63 1.49 4.63 1.37 5.15 1.37 5.15 1.67 5.51 1.67 5.51 0.74 5.57 0.74 5.57 0.62 5.69 0.62 ;
      POLYGON 5.09 1.17 4.51 1.17 4.51 1.73 4.35 1.73 4.35 1.87 4.23 1.87 4.23 1.61 4.39 1.61 4.39 1.17 4.33 1.17 4.33 0.62 4.45 0.62 4.45 1.05 5.09 1.05 ;
      POLYGON 3.97 0.8 3.91 0.8 3.91 1.63 3.93 1.63 3.93 1.87 3.81 1.87 3.81 1.75 3.79 1.75 3.79 1.28 2.95 1.28 2.95 1.16 3.79 1.16 3.79 0.8 3.73 0.8 3.73 0.68 3.97 0.68 ;
      POLYGON 1.14 1.58 1.02 1.58 1.02 1.385 0.99 1.385 0.99 1.2 0.375 1.2 0.375 1.08 0.99 1.08 0.99 0.68 1.11 0.68 1.11 1.265 1.14 1.265 ;
  END
END EDFFTRX1

MACRO DFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX1 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 1.21 2.14 1.33 ;
        RECT 2.02 1.09 2.14 1.33 ;
        RECT 1.81 1.465 1.98 1.725 ;
        RECT 1.86 1.21 1.98 1.725 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.395 1.45 6.655 1.67 ;
        RECT 6.435 1.36 6.555 1.75 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.38 0.68 1.5 2.08 ;
        RECT 1.23 0.885 1.5 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.515 -0.18 6.635 0.76 ;
        RECT 4.955 0.35 5.195 0.47 ;
        RECT 4.955 -0.18 5.075 0.47 ;
        RECT 3.235 -0.18 3.355 0.86 ;
        RECT 1.8 -0.18 1.92 0.73 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 6.495 1.87 6.615 2.79 ;
        RECT 4.895 2.29 5.135 2.79 ;
        RECT 3.115 2.29 3.355 2.79 ;
        RECT 1.86 2.07 1.98 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.175 1.48 7.035 1.48 7.035 1.99 6.915 1.99 6.915 1.36 7.055 1.36 7.055 0.86 6.925 0.86 6.925 1 6.275 1 6.275 0.5 5.435 0.5 5.435 0.71 4.715 0.71 4.715 0.5 4.355 0.5 4.355 1.07 4.435 1.07 4.435 1.31 4.315 1.31 4.315 1.19 3.895 1.19 3.895 1.65 3.775 1.65 3.775 1.07 4.235 1.07 4.235 0.38 4.835 0.38 4.835 0.59 5.315 0.59 5.315 0.38 5.515 0.38 5.515 0.36 5.755 0.36 5.755 0.38 6.395 0.38 6.395 0.88 6.805 0.88 6.805 0.74 6.995 0.74 6.995 0.62 7.115 0.62 7.115 0.74 7.175 0.74 ;
      POLYGON 6.935 1.24 6.275 1.24 6.275 1.34 6.075 1.34 6.075 2.17 2.305 2.17 2.305 1.55 2.28 1.55 2.28 0.68 2.4 0.68 2.4 1.43 2.425 1.43 2.425 2.05 4.175 2.05 4.175 1.67 4.155 1.67 4.155 1.43 4.275 1.43 4.275 1.55 4.295 1.55 4.295 2.05 5.955 2.05 5.955 1.67 5.515 1.67 5.515 1.43 5.635 1.43 5.635 1.55 5.955 1.55 5.955 1.12 6.935 1.12 ;
      POLYGON 5.935 1 5.835 1 5.835 1.31 5.395 1.31 5.395 1.79 5.715 1.79 5.715 1.81 5.835 1.81 5.835 1.93 5.595 1.93 5.595 1.91 5.275 1.91 5.275 1.55 4.915 1.55 4.915 1.67 4.795 1.67 4.795 1.43 5.275 1.43 5.275 1.19 5.715 1.19 5.715 0.88 5.815 0.88 5.815 0.62 5.935 0.62 ;
      POLYGON 5.155 1.29 4.675 1.29 4.675 1.93 4.415 1.93 4.415 1.81 4.555 1.81 4.555 0.95 4.475 0.95 4.475 0.62 4.595 0.62 4.595 0.83 4.675 0.83 4.675 1.17 5.155 1.17 ;
      POLYGON 4.115 0.8 3.655 0.8 3.655 1.77 3.935 1.77 3.935 1.81 4.055 1.81 4.055 1.93 3.815 1.93 3.815 1.89 3.535 1.89 3.535 1.67 2.935 1.67 2.935 1.43 3.055 1.43 3.055 1.55 3.535 1.55 3.535 0.68 4.115 0.68 ;
      POLYGON 3.415 1.43 3.295 1.43 3.295 1.31 2.815 1.31 2.815 1.81 2.875 1.81 2.875 1.93 2.635 1.93 2.635 1.81 2.695 1.81 2.695 0.74 2.795 0.74 2.795 0.56 2.16 0.56 2.16 0.97 1.74 0.97 1.74 1.24 1.62 1.24 1.62 0.85 2.04 0.85 2.04 0.44 2.915 0.44 2.915 0.86 2.815 0.86 2.815 1.19 3.415 1.19 ;
      POLYGON 1.11 1.58 0.99 1.58 0.99 1.2 0.375 1.2 0.375 1.08 0.99 1.08 0.99 0.68 1.11 0.68 ;
  END
END DFFX1

MACRO MDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX8 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.345 2.775 2.19 ;
        RECT 2.655 0.665 2.775 0.985 ;
        RECT 2.635 0.865 2.755 1.465 ;
        RECT 0.07 1.025 2.755 1.145 ;
        RECT 1.815 0.665 1.935 2.19 ;
        RECT 0.975 0.665 1.095 2.185 ;
        RECT 0.135 0.665 0.255 2.185 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 1.155 5.205 1.38 ;
        RECT 5.085 0.98 5.205 1.38 ;
    END
  END CK
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.535 1.2 9.655 1.44 ;
        RECT 9.35 1.2 9.655 1.435 ;
        RECT 9.35 1.175 9.5 1.435 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.745 1.21 11.115 1.395 ;
        RECT 10.745 1.21 11.005 1.42 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.275 0.97 11.395 1.21 ;
        RECT 11.035 0.94 11.295 1.09 ;
        RECT 10.275 0.97 11.395 1.09 ;
        RECT 10.015 1 10.395 1.12 ;
        RECT 10.015 1 10.135 1.44 ;
    END
  END S0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 11.075 -0.18 11.195 0.82 ;
        RECT 9.795 -0.18 9.915 0.64 ;
        RECT 7.425 -0.18 7.665 0.37 ;
        RECT 5.325 -0.18 5.565 0.38 ;
        RECT 3.915 -0.18 4.035 0.65 ;
        RECT 3.075 -0.18 3.195 0.65 ;
        RECT 2.235 -0.18 2.355 0.655 ;
        RECT 1.395 -0.18 1.515 0.655 ;
        RECT 0.555 -0.18 0.675 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 10.915 1.78 11.035 2.79 ;
        RECT 9.535 1.85 9.655 2.79 ;
        RECT 7.425 2.07 7.665 2.19 ;
        RECT 7.425 2.07 7.545 2.79 ;
        RECT 5.645 2.1 5.765 2.79 ;
        RECT 3.975 1.54 4.095 2.79 ;
        RECT 3.075 1.445 3.195 2.79 ;
        RECT 2.235 1.445 2.355 2.79 ;
        RECT 1.395 1.445 1.515 2.79 ;
        RECT 0.555 1.445 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.635 1.68 11.555 1.68 11.555 1.8 11.435 1.8 11.435 1.66 10.415 1.66 10.415 1.24 10.535 1.24 10.535 1.54 11.515 1.54 11.515 0.85 11.495 0.85 11.495 0.58 11.615 0.58 11.615 0.73 11.635 0.73 ;
      POLYGON 10.555 0.85 10.155 0.85 10.155 0.88 9.895 0.88 9.895 1.56 10.295 1.56 10.295 2.21 10.175 2.21 10.175 1.68 8.985 1.68 8.985 1.76 8.745 1.76 8.745 1.53 8.865 1.53 8.865 0.72 8.785 0.72 8.785 0.6 9.025 0.6 9.025 0.72 8.985 0.72 8.985 1.56 9.775 1.56 9.775 0.76 10.035 0.76 10.035 0.73 10.435 0.73 10.435 0.59 10.555 0.59 ;
      POLYGON 9.435 0.83 9.315 0.83 9.315 0.48 8.665 0.48 8.665 1.15 8.705 1.15 8.705 1.39 8.665 1.39 8.665 1.41 8.625 1.41 8.625 1.88 9.175 1.88 9.175 2.03 9.295 2.03 9.295 2.15 9.055 2.15 9.055 2 8.505 2 8.505 1.29 8.545 1.29 8.545 0.48 8.065 0.48 8.065 0.88 8.145 0.88 8.145 1.12 7.945 1.12 7.945 0.61 7.185 0.61 7.185 0.48 6.705 0.48 6.705 0.97 6.965 0.97 6.965 1.21 6.845 1.21 6.845 1.09 6.585 1.09 6.585 0.36 7.305 0.36 7.305 0.49 7.945 0.49 7.945 0.36 9.435 0.36 ;
      POLYGON 8.425 0.72 8.385 0.72 8.385 1.99 8.265 1.99 8.265 1.36 7.465 1.36 7.465 1.31 7.325 1.31 7.325 1.19 7.585 1.19 7.585 1.24 8.265 1.24 8.265 0.72 8.185 0.72 8.185 0.6 8.425 0.6 ;
      POLYGON 8.225 2.25 7.985 2.25 7.985 1.95 7.045 1.95 7.045 2.23 5.925 2.23 5.925 0.86 4.825 0.86 4.825 1.5 5.245 1.5 5.245 1.74 5.125 1.74 5.125 1.62 4.705 1.62 4.705 0.6 4.965 0.6 4.965 0.74 6.045 0.74 6.045 2.11 6.585 2.11 6.585 1.33 6.425 1.33 6.425 1.21 6.705 1.21 6.705 2.11 6.925 2.11 6.925 1.83 8.105 1.83 8.105 2.13 8.225 2.13 ;
      POLYGON 7.825 1.12 7.705 1.12 7.705 1.07 7.205 1.07 7.205 1.45 7.125 1.45 7.125 1.71 7.005 1.71 7.005 1.33 7.085 1.33 7.085 0.85 6.825 0.85 6.825 0.6 7.065 0.6 7.065 0.73 7.205 0.73 7.205 0.95 7.705 0.95 7.705 0.88 7.825 0.88 ;
      POLYGON 6.465 1.99 6.345 1.99 6.345 1.57 6.185 1.57 6.185 0.62 5.085 0.62 5.085 0.48 4.275 0.48 4.275 1.18 4.155 1.18 4.155 0.36 5.205 0.36 5.205 0.5 6.305 0.5 6.305 1.45 6.465 1.45 ;
      POLYGON 5.725 1.98 4.515 1.98 4.515 2.19 4.395 2.19 4.395 1.42 3.675 1.42 3.675 2.19 3.555 2.19 3.555 1.54 3.495 1.54 3.495 1.225 2.875 1.225 2.875 1.105 3.495 1.105 3.495 0.6 3.615 0.6 3.615 1.3 4.395 1.3 4.395 0.6 4.515 0.6 4.515 1.86 5.605 1.86 5.605 1.13 5.725 1.13 ;
  END
END MDFFHQX8

MACRO CLKAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X8 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.115 0.965 3.235 1.235 ;
        RECT 0.595 0.965 3.235 1.085 ;
        RECT 1.595 0.965 1.835 1.115 ;
        RECT 0.415 1.015 0.855 1.135 ;
        RECT 0.595 0.94 0.855 1.135 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.205 2.535 1.325 ;
        RECT 2.045 1.205 2.305 1.38 ;
        RECT 1.295 1.235 2.305 1.355 ;
        RECT 1.175 1.205 1.415 1.325 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.415 1.295 6.535 2.21 ;
        RECT 6.275 0.715 6.515 0.835 ;
        RECT 3.895 1.295 6.535 1.415 ;
        RECT 3.815 0.765 6.395 0.885 ;
        RECT 5.58 1.175 5.73 1.435 ;
        RECT 5.58 0.715 5.7 1.435 ;
        RECT 5.575 1.295 5.695 2.21 ;
        RECT 5.435 0.715 5.7 0.885 ;
        RECT 4.735 1.295 4.855 2.21 ;
        RECT 4.595 0.715 4.835 0.885 ;
        RECT 3.895 1.295 4.015 2.21 ;
        RECT 3.695 0.715 3.935 0.835 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 5.915 -0.18 6.035 0.645 ;
        RECT 5.075 -0.18 5.195 0.645 ;
        RECT 4.175 -0.18 4.295 0.64 ;
        RECT 3.275 0.46 3.515 0.58 ;
        RECT 3.275 -0.18 3.395 0.58 ;
        RECT 1.735 0.485 1.975 0.605 ;
        RECT 1.735 -0.18 1.855 0.605 ;
        RECT 0.315 -0.18 0.435 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 5.995 1.535 6.115 2.79 ;
        RECT 5.155 1.535 5.275 2.79 ;
        RECT 4.315 1.535 4.435 2.79 ;
        RECT 3.415 2.07 3.535 2.79 ;
        RECT 2.695 2.07 2.815 2.79 ;
        RECT 1.855 2.07 1.975 2.79 ;
        RECT 1.015 2.07 1.135 2.79 ;
        RECT 0.135 2.07 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.46 1.175 3.475 1.175 3.475 1.645 0.475 1.645 0.475 1.525 3.355 1.525 3.355 0.845 1.215 0.845 1.215 0.795 1.095 0.795 1.095 0.675 1.335 0.675 1.335 0.725 2.575 0.725 2.575 0.675 2.815 0.675 2.815 0.725 3.475 0.725 3.475 1.055 5.46 1.055 ;
  END
END CLKAND2X8

MACRO OA21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21XL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.595 1.38 0.99 ;
        RECT 1.23 0.595 1.35 1.24 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 1.02 0.89 1.33 ;
        RECT 0.65 1.175 0.8 1.495 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.04 0.51 1.48 ;
        RECT 0.39 0.96 0.51 1.48 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 0.74 2.535 0.86 ;
        RECT 2.1 0.885 2.25 1.145 ;
        RECT 2.13 0.74 2.25 1.145 ;
        RECT 1.85 1.005 2.25 1.125 ;
        RECT 1.85 1.005 1.97 1.72 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.89 -0.18 2.01 0.4 ;
        RECT 0.615 -0.18 0.735 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.43 1.6 1.55 2.79 ;
        RECT 0.29 1.6 0.41 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 1.4 1.62 1.4 1.62 1.48 1.13 1.48 1.13 1.72 1.01 1.72 1.01 1.36 1.5 1.36 1.5 0.66 1.62 0.66 1.62 1.16 1.69 1.16 ;
      POLYGON 1.11 0.9 0.99 0.9 0.99 0.84 0.075 0.84 0.075 0.72 0.99 0.72 0.99 0.66 1.11 0.66 ;
  END
END OA21XL

MACRO OAI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X2 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.065 3.7 1.435 ;
        RECT 3.525 1.01 3.645 1.385 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.18 2.625 1.425 ;
        RECT 2.275 1.18 2.625 1.4 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.04 1.655 1.16 ;
        RECT 0.39 1.04 0.56 1.28 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.28 0.995 1.4 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.28 0.8 1.725 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7616 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.285 0.65 3.645 0.77 ;
        RECT 2.035 0.94 3.405 1.06 ;
        RECT 3.285 0.65 3.405 1.06 ;
        RECT 2.875 1.545 2.995 2.21 ;
        RECT 1.375 1.545 2.995 1.665 ;
        RECT 2.035 0.94 2.155 2.21 ;
        RECT 1.81 1.175 2.155 1.665 ;
        RECT 0.975 1.56 1.495 1.68 ;
        RECT 0.975 1.56 1.095 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 1.755 0.46 1.995 0.58 ;
        RECT 1.755 -0.18 1.875 0.58 ;
        RECT 0.915 0.46 1.155 0.58 ;
        RECT 0.915 -0.18 1.035 0.58 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.295 1.56 3.415 2.79 ;
        RECT 2.455 1.785 2.575 2.79 ;
        RECT 1.615 1.785 1.735 2.79 ;
        RECT 0.335 1.56 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.005 0.65 3.885 0.65 3.885 0.53 3.165 0.53 3.165 0.65 3.045 0.65 3.045 0.53 2.385 0.53 2.385 0.58 2.145 0.58 2.145 0.46 2.265 0.46 2.265 0.41 4.005 0.41 ;
      POLYGON 2.805 0.77 2.685 0.77 2.685 0.82 0.555 0.82 0.555 0.58 0.675 0.58 0.675 0.7 1.395 0.7 1.395 0.58 1.515 0.58 1.515 0.7 2.565 0.7 2.565 0.65 2.805 0.65 ;
  END
END OAI211X2

MACRO TBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.945 0.78 1.185 0.9 ;
        RECT 0.445 0.86 1.065 0.98 ;
        RECT 0.445 0.86 0.565 1.22 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.175 0.98 2.415 1.1 ;
        RECT 1.115 1.76 2.295 1.88 ;
        RECT 2.175 0.98 2.295 1.88 ;
        RECT 0.885 1.67 1.235 1.79 ;
        RECT 0.885 1.52 1.145 1.79 ;
        RECT 0.885 1.1 1.005 1.79 ;
        RECT 0.725 1.1 1.005 1.22 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.095 1.145 3.215 1.88 ;
        RECT 2.97 0.885 3.12 1.265 ;
        RECT 2.935 0.59 3.055 1.025 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.355 -0.18 3.475 0.64 ;
        RECT 2.455 0.5 2.695 0.62 ;
        RECT 2.455 -0.18 2.575 0.62 ;
        RECT 1.675 -0.18 1.795 0.68 ;
        RECT 0.865 -0.18 0.985 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.515 1.34 3.635 2.79 ;
        RECT 2.555 2.24 2.795 2.79 ;
        RECT 0.945 2.24 1.185 2.79 ;
        RECT 0.135 1.58 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.155 2.25 2.915 2.25 2.915 2.12 0.555 2.12 0.555 1.46 0.065 1.46 0.065 0.62 0.225 0.62 0.225 0.4 0.345 0.4 0.345 0.74 0.185 0.74 0.185 1.34 0.675 1.34 0.675 2 3.035 2 3.035 2.13 3.155 2.13 ;
      POLYGON 2.715 1.15 2.595 1.15 2.595 0.86 2.055 0.86 2.055 1.64 1.815 1.64 1.815 1.52 1.935 1.52 1.935 0.74 2.095 0.74 2.095 0.44 2.215 0.44 2.215 0.74 2.715 0.74 ;
      POLYGON 1.815 1.02 1.545 1.02 1.545 1.52 1.665 1.52 1.665 1.64 1.425 1.64 1.425 0.66 1.285 0.66 1.285 0.4 1.405 0.4 1.405 0.54 1.545 0.54 1.545 0.9 1.815 0.9 ;
  END
END TBUFX2

MACRO DFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX4 0 0 ;
  SIZE 14.21 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.065 0.51 1.55 ;
        RECT 0.36 1.065 0.51 1.52 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 1.41 1.265 1.555 ;
        RECT 0.885 1.5 1.145 1.67 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.675 1.12 4.955 1.24 ;
        RECT 4.655 1.23 4.95 1.38 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.2 1.23 5.495 1.38 ;
        RECT 5.215 1.12 5.495 1.38 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.915 0.74 11.115 0.86 ;
        RECT 10.935 1.42 11.055 2.19 ;
        RECT 10.635 1.42 11.055 1.54 ;
        RECT 9.93 1.3 10.755 1.42 ;
        RECT 9.975 0.74 10.095 2.19 ;
        RECT 9.93 1.175 10.095 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.835 0.74 13.035 0.86 ;
        RECT 12.655 1.42 12.775 2.19 ;
        RECT 12.475 1.42 12.775 1.54 ;
        RECT 11.99 1.3 12.595 1.42 ;
        RECT 11.815 1.42 12.11 1.54 ;
        RECT 11.99 0.74 12.11 1.54 ;
        RECT 11.96 0.74 12.11 1.145 ;
        RECT 11.815 1.42 11.935 2.19 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.21 0.18 ;
        RECT 13.395 -0.18 13.515 0.73 ;
        RECT 12.315 -0.18 12.555 0.38 ;
        RECT 11.355 -0.18 11.595 0.38 ;
        RECT 10.395 -0.18 10.635 0.38 ;
        RECT 9.315 0.64 9.555 0.76 ;
        RECT 9.315 -0.18 9.435 0.76 ;
        RECT 8.535 -0.18 8.655 0.86 ;
        RECT 5.035 0.64 5.275 0.76 ;
        RECT 5.155 -0.18 5.275 0.76 ;
        RECT 2.385 -0.18 2.625 0.36 ;
        RECT 0.625 -0.18 0.745 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.21 2.79 ;
        RECT 13.075 1.54 13.195 2.79 ;
        RECT 12.235 1.54 12.355 2.79 ;
        RECT 11.395 1.54 11.515 2.79 ;
        RECT 10.395 1.54 10.515 2.79 ;
        RECT 9.555 1.6 9.675 2.79 ;
        RECT 8.71 1.76 8.83 2.79 ;
        RECT 7.65 1.88 7.77 2.79 ;
        RECT 4.895 1.98 5.015 2.79 ;
        RECT 4.775 1.98 5.015 2.1 ;
        RECT 3.215 2.16 3.335 2.79 ;
        RECT 3.095 2.16 3.335 2.28 ;
        RECT 2.245 2.16 2.485 2.28 ;
        RECT 2.245 2.16 2.365 2.79 ;
        RECT 0.965 1.79 1.085 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.935 0.92 13.775 0.92 13.775 1.42 13.615 1.42 13.615 2.19 13.495 2.19 13.495 1.42 12.895 1.42 12.895 1.28 13.135 1.28 13.135 1.3 13.655 1.3 13.655 0.8 13.815 0.8 13.815 0.68 13.935 0.68 ;
      POLYGON 13.535 1.18 13.295 1.18 13.295 0.97 13.155 0.97 13.155 0.62 9.795 0.62 9.795 1 9.23 1 9.23 1.28 9.81 1.28 9.81 1.4 9.25 1.4 9.25 2.12 9.13 2.12 9.13 1.4 9.11 1.4 9.11 1.14 7.995 1.14 7.995 1.02 8.955 1.02 8.955 0.68 9.075 0.68 9.075 0.88 9.675 0.88 9.675 0.5 13.275 0.5 13.275 0.85 13.415 0.85 13.415 1.06 13.535 1.06 ;
      POLYGON 8.99 1.52 6.525 1.52 6.525 1.89 6.405 1.89 6.405 0.92 6.385 0.92 6.385 0.68 6.505 0.68 6.505 0.8 6.525 0.8 6.525 1.4 8.87 1.4 8.87 1.26 8.99 1.26 ;
      POLYGON 8.47 1.94 8.205 1.94 8.205 1.76 7.53 1.76 7.53 1.81 6.765 1.81 6.765 1.69 7.41 1.69 7.41 1.64 8.325 1.64 8.325 1.82 8.47 1.82 ;
      POLYGON 8.235 0.86 8.115 0.86 8.115 0.5 7.575 0.5 7.575 0.68 7.455 0.68 7.455 0.8 7.215 0.8 7.215 0.68 7.335 0.68 7.335 0.56 7.455 0.56 7.455 0.38 8.235 0.38 ;
      POLYGON 7.815 1.04 6.975 1.04 6.975 0.92 6.885 0.92 6.885 0.68 7.005 0.68 7.005 0.8 7.095 0.8 7.095 0.92 7.695 0.92 7.695 0.62 7.815 0.62 ;
      POLYGON 7.615 1.28 6.735 1.28 6.735 1.16 6.645 1.16 6.645 0.56 5.705 0.56 5.705 0.74 5.735 0.74 5.735 1.62 5.615 1.62 5.615 1 4.795 1 4.795 0.5 4.38 0.5 4.38 0.48 3.995 0.48 3.995 0.36 4.5 0.36 4.5 0.38 4.915 0.38 4.915 0.88 5.575 0.88 5.575 0.62 5.585 0.62 5.585 0.44 6.765 0.44 6.765 1.04 6.855 1.04 6.855 1.16 7.615 1.16 ;
      POLYGON 6.785 2.25 5.665 2.25 5.665 2.13 5.135 2.13 5.135 1.86 4.055 1.86 4.055 1.56 2.725 1.56 2.725 1.44 2.845 1.44 2.845 0.94 2.005 0.94 2.005 1.22 1.885 1.22 1.885 0.82 2.845 0.82 2.845 0.72 3.105 0.72 3.105 0.84 2.965 0.84 2.965 1.44 4.175 1.44 4.175 1.74 5.255 1.74 5.255 2.01 5.785 2.01 5.785 2.13 6.165 2.13 6.165 1.28 6.125 1.28 6.125 1.04 6.285 1.04 6.285 2.13 6.785 2.13 ;
      POLYGON 6.085 0.92 6.005 0.92 6.005 1.77 6.045 1.77 6.045 2.01 5.925 2.01 5.925 1.89 5.375 1.89 5.375 1.62 4.295 1.62 4.295 1.5 4.415 1.5 4.415 1.32 3.275 1.32 3.275 0.5 3.06 0.5 3.06 0.6 2.145 0.6 2.145 0.52 2.025 0.52 2.025 0.4 2.265 0.4 2.265 0.48 2.94 0.48 2.94 0.38 3.875 0.38 3.875 0.68 4.315 0.68 4.315 0.8 3.755 0.8 3.755 0.5 3.395 0.5 3.395 1.2 4.535 1.2 4.535 1.5 5.495 1.5 5.495 1.77 5.885 1.77 5.885 0.8 5.965 0.8 5.965 0.68 6.085 0.68 ;
      POLYGON 4.675 1 4.555 1 4.555 1.04 3.515 1.04 3.515 0.62 3.635 0.62 3.635 0.92 4.435 0.92 4.435 0.88 4.555 0.88 4.555 0.62 4.675 0.62 ;
      POLYGON 4.655 2.25 4.08 2.25 4.08 2.1 3.815 2.1 3.815 1.8 2.485 1.8 2.485 1.48 1.645 1.48 1.645 0.54 1.285 0.54 1.285 1.24 1.165 1.24 1.165 0.945 0.24 0.945 0.24 1.67 0.585 1.67 0.585 1.91 0.465 1.91 0.465 1.79 0.12 1.79 0.12 0.78 0.145 0.78 0.145 0.66 0.265 0.66 0.265 0.825 1.165 0.825 1.165 0.42 1.765 0.42 1.765 1.36 2.485 1.36 2.485 1.06 2.625 1.06 2.625 1.3 2.605 1.3 2.605 1.68 3.935 1.68 3.935 1.98 4.2 1.98 4.2 2.13 4.655 2.13 ;
      POLYGON 3.695 2.16 3.455 2.16 3.455 2.04 1.605 2.04 1.605 1.8 1.405 1.8 1.405 0.66 1.525 0.66 1.525 1.68 1.725 1.68 1.725 1.92 3.575 1.92 3.575 2.04 3.695 2.04 ;
  END
END DFFSRX4

MACRO ADDHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.52 0.36 2.8 0.48 ;
        RECT 2.04 0.65 2.64 0.77 ;
        RECT 2.52 0.36 2.64 0.77 ;
        RECT 2.04 0.38 2.16 0.77 ;
        RECT 0.89 0.38 2.16 0.5 ;
        RECT 0.735 0.71 1.01 0.83 ;
        RECT 0.89 0.38 1.01 0.83 ;
        RECT 0.73 0.98 0.97 1.1 ;
        RECT 0.595 0.94 0.855 1.09 ;
        RECT 0.735 0.71 0.855 1.1 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.14 0.9 1.435 1.135 ;
        RECT 1.13 0.9 1.435 1.11 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 0.6 0.29 2.21 ;
        RECT 0.07 1.175 0.29 1.435 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.38 1.175 4.57 1.435 ;
        RECT 4.38 0.8 4.5 1.435 ;
        RECT 4.36 1.3 4.48 1.99 ;
        RECT 4.36 0.68 4.48 0.92 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.88 0.68 4.12 0.8 ;
        RECT 3.98 -0.18 4.1 0.8 ;
        RECT 2.28 -0.18 2.4 0.53 ;
        RECT 0.53 0.47 0.77 0.59 ;
        RECT 0.65 -0.18 0.77 0.59 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.94 1.72 4.06 2.79 ;
        RECT 2.22 1.85 2.46 1.97 ;
        RECT 2.22 1.85 2.34 2.79 ;
        RECT 1.49 2.02 1.61 2.79 ;
        RECT 0.53 1.91 0.77 2.15 ;
        RECT 0.53 1.91 0.65 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.26 1.18 4.02 1.18 4.02 1.12 3.88 1.12 3.88 1.6 3.42 1.6 3.42 1.87 3.3 1.87 3.3 1.48 3.76 1.48 3.76 1.12 3.3 1.12 3.3 0.86 3.18 0.86 3.18 0.62 3.3 0.62 3.3 0.74 3.42 0.74 3.42 1 4.14 1 4.14 1.06 4.26 1.06 ;
      POLYGON 3.86 0.48 3.74 0.48 3.74 0.5 3.04 0.5 3.04 0.74 2.88 0.74 2.88 1.01 2.74 1.01 2.74 1.37 2.94 1.37 2.94 1.87 2.82 1.87 2.82 1.49 2.62 1.49 2.62 0.89 2.76 0.89 2.76 0.62 2.92 0.62 2.92 0.38 3.62 0.38 3.62 0.36 3.86 0.36 ;
      POLYGON 3.64 1.36 3.18 1.36 3.18 2.11 2.58 2.11 2.58 1.73 1.92 1.73 1.92 1.87 1.8 1.87 1.8 0.62 1.92 0.62 1.92 1.61 2.7 1.61 2.7 1.99 3.06 1.99 3.06 1.25 2.86 1.25 2.86 1.13 3.18 1.13 3.18 1.24 3.64 1.24 ;
      POLYGON 1.675 1.375 1.13 1.375 1.13 2.09 1.01 2.09 1.01 1.375 0.57 1.375 0.57 1.48 0.45 1.48 0.45 1.24 0.57 1.24 0.57 1.255 1.555 1.255 1.555 0.78 1.23 0.78 1.23 0.66 1.675 0.66 ;
  END
END ADDHX1

MACRO EDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFXL 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.13 0.51 1.6 ;
        RECT 0.38 1.13 0.5 1.63 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.39 1.195 6.655 1.445 ;
        RECT 6.395 1.175 6.655 1.445 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.03 1.175 7.18 1.435 ;
        RECT 6.89 1.195 7.18 1.435 ;
        RECT 5.77 1.565 6.97 1.685 ;
        RECT 6.85 1.315 6.97 1.685 ;
        RECT 5.27 2.13 5.89 2.25 ;
        RECT 5.77 0.96 5.89 2.25 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.54 0.74 7.78 0.86 ;
        RECT 7.61 0.74 7.76 1.145 ;
        RECT 7.6 1.005 7.72 1.58 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.315 0.68 9.435 2.09 ;
        RECT 9.06 1.465 9.435 1.725 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.895 -0.18 9.015 0.92 ;
        RECT 8.08 -0.18 8.2 0.4 ;
        RECT 6.61 0.455 6.85 0.575 ;
        RECT 6.61 -0.18 6.73 0.575 ;
        RECT 4.59 0.68 4.83 0.8 ;
        RECT 4.59 -0.18 4.71 0.8 ;
        RECT 2.57 0.6 2.81 0.72 ;
        RECT 2.57 -0.18 2.69 0.72 ;
        RECT 0.56 -0.18 0.68 0.77 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.895 1.97 9.015 2.79 ;
        RECT 8.08 1.98 8.2 2.79 ;
        RECT 6.61 1.805 6.85 1.925 ;
        RECT 6.61 1.805 6.73 2.79 ;
        RECT 4.59 2.23 4.71 2.79 ;
        RECT 2.69 2.04 2.81 2.79 ;
        RECT 2.57 2.04 2.81 2.16 ;
        RECT 0.56 1.75 0.68 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.195 1.34 8.68 1.34 8.68 1.58 8.56 1.58 8.56 0.92 8.505 0.92 8.505 0.68 8.625 0.68 8.625 0.8 8.68 0.8 8.68 1.22 9.195 1.22 ;
      POLYGON 7.94 0.52 7.45 0.52 7.45 0.5 7.09 0.5 7.09 0.815 6.175 0.815 6.175 0.5 5.19 0.5 5.19 0.86 5.17 0.86 5.17 1.65 5.25 1.65 5.25 1.77 5.01 1.77 5.01 1.65 5.05 1.65 5.05 1.49 4.43 1.49 4.43 1.25 4.55 1.25 4.55 1.37 5.05 1.37 5.05 0.74 5.07 0.74 5.07 0.38 6.295 0.38 6.295 0.695 6.97 0.695 6.97 0.38 7.57 0.38 7.57 0.4 7.94 0.4 ;
      POLYGON 7.42 1.77 7.09 1.77 7.09 1.65 7.3 1.65 7.3 1.055 6.23 1.055 6.23 1.44 6.11 1.44 6.11 0.935 7.21 0.935 7.21 0.62 7.33 0.62 7.33 0.815 7.42 0.815 ;
      POLYGON 5.65 2.01 4.3 2.01 4.3 2.09 3.65 2.09 3.65 2.01 3.17 2.01 3.17 1.68 2.21 1.68 2.21 2.01 1.49 2.01 1.49 1.95 1.37 1.95 1.37 0.62 1.49 0.62 1.49 1.83 1.61 1.83 1.61 1.89 2.09 1.89 2.09 1.56 3.29 1.56 3.29 1.89 3.77 1.89 3.77 1.97 4.18 1.97 4.18 1.89 5.53 1.89 5.53 0.62 5.65 0.62 ;
      POLYGON 4.93 1.25 4.81 1.25 4.81 1.13 4.31 1.13 4.31 1.73 4.01 1.73 4.01 1.85 3.89 1.85 3.89 1.61 4.19 1.61 4.19 1.13 3.89 1.13 3.89 0.62 4.01 0.62 4.01 1.01 4.93 1.01 ;
      POLYGON 4.07 1.49 3.95 1.49 3.95 1.37 3.65 1.37 3.65 1.2 3.41 1.2 3.41 0.96 3.65 0.96 3.65 0.56 3.05 0.56 3.05 0.96 2.33 0.96 2.33 0.5 1.73 0.5 1.73 1.49 1.61 1.49 1.61 0.5 1.1 0.5 1.1 1.87 0.98 1.87 0.98 0.38 2.01 0.38 2.01 0.36 2.25 0.36 2.25 0.38 2.45 0.38 2.45 0.84 2.93 0.84 2.93 0.44 3.77 0.44 3.77 1.25 4.07 1.25 ;
      POLYGON 3.65 1.77 3.41 1.77 3.41 1.44 2.37 1.44 2.37 1.32 3.17 1.32 3.17 0.68 3.41 0.68 3.41 0.8 3.29 0.8 3.29 1.32 3.53 1.32 3.53 1.65 3.65 1.65 ;
      POLYGON 3.53 2.25 2.93 2.25 2.93 1.92 2.45 1.92 2.45 2.25 1.99 2.25 1.99 2.13 2.33 2.13 2.33 1.8 3.05 1.8 3.05 2.13 3.53 2.13 ;
      POLYGON 3.03 1.2 1.97 1.2 1.97 1.77 1.73 1.77 1.73 1.65 1.85 1.65 1.85 0.68 2.09 0.68 2.09 0.8 1.97 0.8 1.97 1.08 3.03 1.08 ;
      POLYGON 0.84 1.13 0.72 1.13 0.72 1.01 0.24 1.01 0.24 1.72 0.26 1.72 0.26 1.96 0.14 1.96 0.14 1.84 0.12 1.84 0.12 0.77 0.14 0.77 0.14 0.53 0.26 0.53 0.26 0.89 0.84 0.89 ;
  END
END EDFFXL

MACRO CLKINVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX20 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.16 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.165 6.365 1.285 ;
        RECT 0.885 1.165 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.285 1.45 7.405 2.21 ;
        RECT 0.555 0.925 7.405 1.045 ;
        RECT 7.285 0.4 7.405 1.045 ;
        RECT 0.565 1.5 7.405 1.62 ;
        RECT 6.74 1.175 6.89 1.62 ;
        RECT 6.485 1.315 6.89 1.62 ;
        RECT 6.485 0.925 6.605 1.62 ;
        RECT 6.445 1.445 6.565 2.21 ;
        RECT 6.445 0.4 6.565 1.045 ;
        RECT 5.605 1.445 5.725 2.21 ;
        RECT 5.605 0.4 5.725 1.045 ;
        RECT 4.765 1.445 4.885 2.21 ;
        RECT 4.765 0.4 4.885 1.045 ;
        RECT 3.925 1.445 4.045 2.21 ;
        RECT 3.925 0.4 4.045 1.045 ;
        RECT 3.085 1.445 3.205 2.21 ;
        RECT 3.085 0.4 3.205 1.045 ;
        RECT 2.245 1.445 2.365 2.21 ;
        RECT 2.245 0.4 2.365 1.045 ;
        RECT 1.405 1.445 1.525 2.21 ;
        RECT 1.395 0.4 1.515 1.045 ;
        RECT 0.565 1.445 0.685 2.21 ;
        RECT 0.555 0.4 0.675 1.045 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.865 -0.18 6.985 0.805 ;
        RECT 6.025 -0.18 6.145 0.805 ;
        RECT 5.185 -0.18 5.305 0.805 ;
        RECT 4.345 -0.18 4.465 0.805 ;
        RECT 3.505 -0.18 3.625 0.805 ;
        RECT 2.665 -0.18 2.785 0.805 ;
        RECT 1.825 -0.18 1.945 0.805 ;
        RECT 0.975 -0.18 1.095 0.805 ;
        RECT 0.135 -0.18 0.255 0.91 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.865 1.74 6.985 2.79 ;
        RECT 6.025 1.74 6.145 2.79 ;
        RECT 5.185 1.74 5.305 2.79 ;
        RECT 4.345 1.74 4.465 2.79 ;
        RECT 3.505 1.74 3.625 2.79 ;
        RECT 2.665 1.74 2.785 2.79 ;
        RECT 1.825 1.74 1.945 2.79 ;
        RECT 0.985 1.74 1.105 2.79 ;
        RECT 0.145 1.445 0.265 2.79 ;
    END
  END VDD
END CLKINVX20

MACRO MX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X8 0 0 ;
  SIZE 5.8 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.12 1.505 1.24 ;
        RECT 0.645 1.5 1.385 1.62 ;
        RECT 1.265 1.12 1.385 1.62 ;
        RECT 0.645 1.175 0.765 1.62 ;
        RECT 0.36 1.175 0.765 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.11 1.145 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.08 2.54 1.46 ;
        RECT 2.28 1.08 2.54 1.275 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.725 0.765 5.465 0.885 ;
        RECT 5.345 0.645 5.465 0.885 ;
        RECT 5.34 0.765 5.46 2.205 ;
        RECT 2.97 1.225 5.46 1.345 ;
        RECT 4.445 0.715 4.685 0.885 ;
        RECT 4.5 1.225 4.62 2.205 ;
        RECT 3.605 0.715 3.845 0.835 ;
        RECT 3.66 1.225 3.78 2.21 ;
        RECT 2.97 1.175 3.12 1.435 ;
        RECT 2.82 1.345 3.09 1.465 ;
        RECT 2.97 0.6 3.09 1.465 ;
        RECT 2.765 0.6 3.09 0.72 ;
        RECT 2.82 1.345 2.94 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.8 0.18 ;
        RECT 4.925 -0.18 5.045 0.645 ;
        RECT 4.085 -0.18 4.205 0.645 ;
        RECT 3.245 -0.18 3.365 0.645 ;
        RECT 2.345 0.46 2.585 0.58 ;
        RECT 2.345 -0.18 2.465 0.58 ;
        RECT 0.825 -0.18 0.945 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.8 2.79 ;
        RECT 4.92 1.465 5.04 2.79 ;
        RECT 4.08 1.465 4.2 2.79 ;
        RECT 3.24 1.465 3.36 2.79 ;
        RECT 2.4 1.58 2.52 2.79 ;
        RECT 0.96 1.74 1.2 2.14 ;
        RECT 0.96 1.74 1.08 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.8 1.215 2.68 1.215 2.68 0.96 2.16 0.96 2.16 1.78 1.78 1.78 1.78 2.2 1.66 2.2 1.66 1.66 2.04 1.66 2.04 0.96 1.985 0.96 1.985 0.75 1.765 0.75 1.765 0.5 1.885 0.5 1.885 0.63 2.105 0.63 2.105 0.84 2.8 0.84 ;
      POLYGON 1.92 1.54 1.625 1.54 1.625 0.99 0.24 0.99 0.24 1.555 0.525 1.555 0.525 1.92 0.405 1.92 0.405 1.675 0.12 1.675 0.12 0.75 0.345 0.75 0.345 0.5 0.465 0.5 0.465 0.87 1.745 0.87 1.745 0.88 1.865 0.88 1.865 1 1.745 1 1.745 1.42 1.92 1.42 ;
  END
END MX2X8

MACRO CLKMX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X6 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 1.555 1.17 1.675 ;
        RECT 1.05 1.35 1.17 1.675 ;
        RECT 0.41 1.195 0.53 1.675 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.045 0.85 1.435 ;
        RECT 0.73 1.035 0.85 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 1.215 2.25 1.435 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.87 1.215 1.99 1.455 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.21 1.43 4.33 2.21 ;
        RECT 3.99 0.8 4.29 0.92 ;
        RECT 4.17 0.405 4.29 0.92 ;
        RECT 4.03 1.43 4.33 1.55 ;
        RECT 4.03 1.19 4.15 1.55 ;
        RECT 3.33 1.04 4.11 1.31 ;
        RECT 3.99 0.8 4.11 1.31 ;
        RECT 3.37 1.04 3.49 2.21 ;
        RECT 3.33 0.405 3.45 1.31 ;
        RECT 2.67 1.19 4.15 1.31 ;
        RECT 2.67 1.175 2.83 1.435 ;
        RECT 2.53 1.36 2.79 1.48 ;
        RECT 2.67 0.63 2.79 1.48 ;
        RECT 2.43 0.63 2.79 0.75 ;
        RECT 2.53 1.36 2.65 2.21 ;
        RECT 2.43 0.4 2.55 0.75 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.75 -0.18 3.87 0.92 ;
        RECT 2.91 -0.18 3.03 0.92 ;
        RECT 2.01 -0.18 2.13 0.74 ;
        RECT 0.73 -0.18 0.85 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.79 1.43 3.91 2.79 ;
        RECT 2.95 1.43 3.07 2.79 ;
        RECT 2.11 1.555 2.23 2.79 ;
        RECT 0.57 1.795 0.69 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.49 1.24 2.37 1.24 2.37 0.99 1.75 0.99 1.75 1.84 1.43 1.84 1.43 2.21 1.31 2.21 1.31 1.72 1.63 1.72 1.63 0.99 1.47 0.99 1.47 0.675 1.37 0.675 1.37 0.435 1.49 0.435 1.49 0.555 1.59 0.555 1.59 0.87 2.49 0.87 ;
      POLYGON 1.51 1.6 1.39 1.6 1.39 1.23 1.23 1.23 1.23 0.915 0.24 0.915 0.24 1.555 0.27 1.555 0.27 2.035 0.15 2.035 0.15 1.675 0.12 1.675 0.12 0.675 0.25 0.675 0.25 0.5 0.37 0.5 0.37 0.795 1.35 0.795 1.35 1.11 1.51 1.11 ;
  END
END CLKMX2X6

MACRO EDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX4 0 0 ;
  SIZE 15.08 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.645 1.41 ;
        RECT 0.525 1.17 0.645 1.41 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 1.25 2.395 1.37 ;
        RECT 1.025 1.81 2.135 1.93 ;
        RECT 2.015 1.25 2.135 1.93 ;
        RECT 1.025 1.17 1.145 1.93 ;
        RECT 0.885 1.52 1.145 1.67 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.655 1.23 5.035 1.42 ;
        RECT 4.655 1.23 4.915 1.445 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.22 9.555 1.45 ;
        RECT 9.305 1.04 9.425 1.45 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.885 1.49 12.125 1.61 ;
        RECT 11.325 0.85 12.105 0.97 ;
        RECT 11.985 0.68 12.105 0.97 ;
        RECT 11.325 1.37 12.005 1.49 ;
        RECT 11.325 1.175 11.53 1.49 ;
        RECT 10.925 1.49 11.445 1.61 ;
        RECT 11.325 0.8 11.445 1.61 ;
        RECT 11.145 0.8 11.445 0.92 ;
        RECT 11.145 0.68 11.265 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.805 1.49 14.045 1.61 ;
        RECT 12.845 1.38 13.925 1.5 ;
        RECT 12.86 0.85 13.785 0.97 ;
        RECT 13.665 0.68 13.785 0.97 ;
        RECT 12.845 1.38 13.085 1.61 ;
        RECT 12.83 1.175 12.98 1.435 ;
        RECT 12.86 0.8 12.98 1.61 ;
        RECT 12.825 0.68 12.945 0.92 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 15.08 0.18 ;
        RECT 14.085 -0.18 14.205 0.73 ;
        RECT 13.245 -0.18 13.365 0.73 ;
        RECT 12.405 -0.18 12.525 0.73 ;
        RECT 11.565 -0.18 11.685 0.73 ;
        RECT 10.725 -0.18 10.845 0.73 ;
        RECT 9.825 -0.18 9.945 0.82 ;
        RECT 8.175 0.7 8.415 0.82 ;
        RECT 8.175 -0.18 8.295 0.82 ;
        RECT 6.455 0.53 6.695 0.65 ;
        RECT 6.455 -0.18 6.575 0.65 ;
        RECT 4.735 -0.18 4.975 0.34 ;
        RECT 3.775 -0.18 3.895 0.38 ;
        RECT 2.645 0.53 2.885 0.65 ;
        RECT 2.645 -0.18 2.765 0.65 ;
        RECT 2.255 0.53 2.495 0.65 ;
        RECT 2.375 -0.18 2.495 0.65 ;
        RECT 0.805 -0.18 0.925 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 15.08 2.79 ;
        RECT 14.285 1.97 14.525 2.09 ;
        RECT 14.285 1.97 14.405 2.79 ;
        RECT 13.325 1.97 13.565 2.09 ;
        RECT 13.325 1.97 13.445 2.79 ;
        RECT 12.365 1.97 12.605 2.09 ;
        RECT 12.365 1.97 12.485 2.79 ;
        RECT 11.405 1.97 11.645 2.09 ;
        RECT 11.405 1.97 11.525 2.79 ;
        RECT 10.445 1.97 10.685 2.09 ;
        RECT 10.445 1.97 10.565 2.79 ;
        RECT 9.565 2.29 9.805 2.79 ;
        RECT 8.335 2.29 8.575 2.79 ;
        RECT 6.555 2.11 6.675 2.79 ;
        RECT 5.255 2.15 5.375 2.79 ;
        RECT 4.445 2.17 4.565 2.79 ;
        RECT 0.785 2.29 1.025 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.945 2.08 14.825 2.08 14.825 1.55 14.585 1.55 14.585 0.97 14.045 0.97 14.045 1.26 13.925 1.26 13.925 0.85 14.505 0.85 14.505 0.68 14.625 0.68 14.625 0.8 14.705 0.8 14.705 1.43 14.945 1.43 ;
      POLYGON 14.465 1.85 10.145 1.85 10.145 1.95 10.04 1.95 10.04 2.17 8.065 2.17 8.065 2.15 7.005 2.15 7.005 1.99 6.33 1.99 6.33 2.03 5.005 2.03 5.005 2.05 3.945 2.05 3.945 2.25 3.825 2.25 3.825 1.93 4.885 1.93 4.885 1.91 6.21 1.91 6.21 1.87 7.125 1.87 7.125 2.03 8.255 2.03 8.255 2.05 9.92 2.05 9.92 1.83 10.025 1.83 10.025 1.43 10.245 1.43 10.245 0.68 10.365 0.68 10.365 1.17 11.045 1.17 11.045 1.29 10.365 1.29 10.365 1.55 10.145 1.55 10.145 1.73 14.345 1.73 14.345 1.09 14.465 1.09 ;
      POLYGON 10.105 1.31 9.905 1.31 9.905 1.71 9.64 1.71 9.64 1.93 8.375 1.93 8.375 1.91 7.455 1.91 7.455 1.55 7.535 1.55 7.535 0.64 7.655 0.64 7.655 1.67 7.575 1.67 7.575 1.79 8.495 1.79 8.495 1.81 9.52 1.81 9.52 1.59 9.785 1.59 9.785 1.19 9.985 1.19 9.985 1.07 10.105 1.07 ;
      POLYGON 9.465 0.92 9.175 0.92 9.175 1.57 9.325 1.57 9.325 1.69 9.055 1.69 9.055 0.8 9.345 0.8 9.345 0.68 9.08 0.68 9.08 0.52 8.655 0.52 8.655 1.06 7.935 1.06 7.935 0.52 7.415 0.52 7.415 1.43 7.295 1.43 7.295 0.52 6.935 0.52 6.935 0.89 6.055 0.89 6.055 1.43 5.935 1.43 5.935 0.48 5.455 0.48 5.455 0.36 6.055 0.36 6.055 0.77 6.815 0.77 6.815 0.4 7.695 0.4 7.695 0.36 7.935 0.36 7.935 0.4 8.055 0.4 8.055 0.94 8.535 0.94 8.535 0.48 8.435 0.48 8.435 0.36 8.675 0.36 8.675 0.4 9.2 0.4 9.2 0.56 9.465 0.56 ;
      POLYGON 8.935 1.69 8.695 1.69 8.695 1.57 8.775 1.57 8.775 1.37 7.775 1.37 7.775 1.25 8.775 1.25 8.775 0.64 8.895 0.64 8.895 1.57 8.935 1.57 ;
      POLYGON 7.175 1.49 7.155 1.49 7.155 1.75 7.035 1.75 7.035 1.49 6.575 1.49 6.575 1.37 6.415 1.37 6.415 1.25 6.695 1.25 6.695 1.37 7.055 1.37 7.055 0.64 7.175 0.64 ;
      POLYGON 6.935 1.25 6.815 1.25 6.815 1.13 6.295 1.13 6.295 1.67 6.035 1.67 6.035 1.69 5.695 1.69 5.695 0.82 5.575 0.82 5.575 0.7 5.815 0.7 5.815 1.55 6.175 1.55 6.175 1.01 6.935 1.01 ;
      POLYGON 5.335 0.48 5.215 0.48 5.215 0.58 4.135 0.58 4.135 0.66 3.685 0.66 3.685 1.13 2.855 1.13 2.855 1.75 2.735 1.75 2.735 1.13 1.825 1.13 1.825 1.57 1.895 1.57 1.895 1.69 1.655 1.69 1.655 1.57 1.705 1.57 1.705 0.72 1.555 0.72 1.555 0.6 1.825 0.6 1.825 1.01 3.565 1.01 3.565 0.54 4.015 0.54 4.015 0.46 5.095 0.46 5.095 0.36 5.335 0.36 ;
      POLYGON 4.955 1.69 4.375 1.69 4.375 1.23 4.175 1.23 4.175 1.11 4.375 1.11 4.375 0.82 4.255 0.82 4.255 0.7 4.495 0.7 4.495 1.57 4.955 1.57 ;
      POLYGON 4.085 1.81 3.965 1.81 3.965 1.57 3.245 1.57 3.245 1.81 3.125 1.81 3.125 1.45 4.085 1.45 ;
      POLYGON 3.665 2.05 2.375 2.05 2.375 1.81 2.255 1.81 2.255 1.69 2.495 1.69 2.495 1.93 3.545 1.93 3.545 1.69 3.665 1.69 ;
      POLYGON 3.245 0.52 3.125 0.52 3.125 0.89 1.945 0.89 1.945 0.48 1.345 0.48 1.345 0.8 1.385 0.8 1.385 1.57 1.505 1.57 1.505 1.69 1.265 1.69 1.265 0.92 1.225 0.92 1.225 0.36 2.065 0.36 2.065 0.77 3.005 0.77 3.005 0.4 3.245 0.4 ;
      POLYGON 2.055 2.17 0.365 2.17 0.365 1.675 0.12 1.675 0.12 0.93 0.385 0.93 0.385 0.68 0.505 0.68 0.505 1.05 0.24 1.05 0.24 1.555 0.485 1.555 0.485 2.05 2.055 2.05 ;
  END
END EDFFTRX4

MACRO NOR2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1 0.51 1.475 ;
        RECT 0.36 1 0.51 1.45 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 1.165 1.255 1.44 ;
        RECT 0.885 1.215 1.255 1.38 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3196 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.59 0.675 0.85 ;
        RECT 0.12 0.76 0.595 0.88 ;
        RECT 0.475 0.73 0.675 0.85 ;
        RECT 0.275 1.595 0.395 2.21 ;
        RECT 0.12 1.595 0.395 1.715 ;
        RECT 0.12 0.76 0.24 1.715 ;
        RECT 0.07 0.885 0.24 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.805 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.915 1.56 1.035 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.8 1.395 1.8 1.395 1.045 1.015 1.045 1.015 1.09 0.715 1.09 0.715 0.97 0.895 0.97 0.895 0.925 1.395 0.925 1.395 0.565 1.515 0.565 ;
  END
END NOR2BX1

MACRO SDFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX1 0 0 ;
  SIZE 12.76 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.27 2.25 1.725 ;
        RECT 2.105 1.25 2.225 1.725 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.885 2.11 7.765 2.23 ;
        RECT 6.885 1.79 7.005 2.23 ;
        RECT 5.245 1.79 7.005 1.91 ;
        RECT 5.245 1.4 5.365 1.91 ;
        RECT 3.515 1.4 5.365 1.52 ;
        RECT 3.515 1.23 3.755 1.52 ;
        RECT 3.395 1.26 3.755 1.38 ;
        RECT 3.495 1.23 3.755 1.38 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.015 1.5 10.365 1.63 ;
        RECT 9.875 1.505 10.135 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.165 1.26 10.705 1.38 ;
        RECT 10.165 1.23 10.425 1.38 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.585 1.27 12.045 1.39 ;
        RECT 11.61 1.23 12.045 1.39 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.165 0.99 12.285 1.23 ;
        RECT 11.905 0.94 12.165 1.11 ;
        RECT 11.065 0.99 12.285 1.11 ;
        RECT 11.605 0.87 11.725 1.11 ;
        RECT 11.065 0.99 11.185 1.63 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 1.32 1.545 2.085 ;
        RECT 1.365 0.65 1.485 0.89 ;
        RECT 1.325 0.77 1.445 1.44 ;
        RECT 1.23 0.885 1.445 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.76 0.18 ;
        RECT 12.085 -0.18 12.205 0.75 ;
        RECT 10.685 0.51 10.925 0.63 ;
        RECT 10.805 -0.18 10.925 0.63 ;
        RECT 9.695 -0.18 9.935 0.32 ;
        RECT 7.825 -0.18 7.945 0.86 ;
        RECT 3.075 -0.18 3.315 0.32 ;
        RECT 1.785 -0.18 1.905 0.89 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.76 2.79 ;
        RECT 11.905 1.93 12.025 2.79 ;
        RECT 10.525 1.99 10.765 2.11 ;
        RECT 10.525 1.99 10.645 2.79 ;
        RECT 9.715 2.29 9.955 2.79 ;
        RECT 7.905 2.23 8.025 2.79 ;
        RECT 6.185 2.29 6.425 2.79 ;
        RECT 4.395 2.12 4.635 2.24 ;
        RECT 4.395 2.12 4.515 2.79 ;
        RECT 3.135 2.12 3.255 2.79 ;
        RECT 1.845 1.725 1.965 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.685 0.69 12.525 0.69 12.525 1.75 12.445 1.75 12.445 2.05 12.325 2.05 12.325 1.63 11.345 1.63 11.345 1.51 12.405 1.51 12.405 0.57 12.685 0.57 ;
      POLYGON 11.565 0.75 11.485 0.75 11.485 0.87 10.945 0.87 10.945 1.75 11.345 1.75 11.345 2.05 11.225 2.05 11.225 1.87 10.825 1.87 10.825 0.87 10.445 0.87 10.445 0.56 9.005 0.56 9.005 0.74 9.025 0.74 9.025 1.82 8.905 1.82 8.905 0.86 8.885 0.86 8.885 0.44 10.565 0.44 10.565 0.75 11.365 0.75 11.365 0.63 11.445 0.63 11.445 0.51 11.565 0.51 ;
      POLYGON 10.325 0.8 10.045 0.8 10.045 1.2 9.755 1.2 9.755 2.05 10.165 2.05 10.165 1.84 10.285 1.84 10.285 2.17 8.525 2.17 8.525 2.2 8.285 2.2 8.285 2 7.885 2 7.885 1.99 7.125 1.99 7.125 1.67 6.745 1.67 6.745 1.41 6.565 1.41 6.565 1.29 6.865 1.29 6.865 1.55 7.245 1.55 7.245 1.87 8.005 1.87 8.005 1.88 8.43 1.88 8.43 2.05 9.635 2.05 9.635 1.2 9.535 1.2 9.535 0.96 9.655 0.96 9.655 1.08 9.925 1.08 9.925 0.68 10.325 0.68 ;
      POLYGON 9.475 1.93 9.235 1.93 9.235 1.5 9.145 1.5 9.145 1.26 9.235 1.26 9.235 0.8 9.215 0.8 9.215 0.68 9.455 0.68 9.455 0.8 9.355 0.8 9.355 1.81 9.475 1.81 ;
      POLYGON 8.665 1.76 8.425 1.76 8.425 1.64 8.465 1.64 8.465 1.19 7.225 1.19 7.225 1.07 8.465 1.07 8.465 0.62 8.585 0.62 8.585 1.64 8.665 1.64 ;
      POLYGON 8.145 1.43 7.485 1.43 7.485 1.63 7.605 1.63 7.605 1.75 7.365 1.75 7.365 1.43 6.985 1.43 6.985 1.17 6.445 1.17 6.445 1.64 5.905 1.64 5.905 1.52 6.325 1.52 6.325 1.08 6.005 1.08 6.005 0.62 6.125 0.62 6.125 0.96 6.445 0.96 6.445 1.05 6.985 1.05 6.985 0.62 7.105 0.62 7.105 1.31 8.145 1.31 ;
      POLYGON 7.525 0.86 7.405 0.86 7.405 0.62 7.225 0.62 7.225 0.5 6.745 0.5 6.745 0.8 6.505 0.8 6.505 0.68 6.625 0.68 6.625 0.38 7.345 0.38 7.345 0.5 7.525 0.5 ;
      POLYGON 6.765 2.17 4.91 2.17 4.91 2 4.235 2 4.235 2.25 4.115 2.25 4.115 2 3.015 2 3.015 2.05 2.385 2.05 2.385 2.085 2.265 2.085 2.265 1.845 2.37 1.845 2.37 1.13 2.265 1.13 2.265 0.65 2.385 0.65 2.385 1.01 2.49 1.01 2.49 1.93 2.895 1.93 2.895 1.88 5.03 1.88 5.03 2.05 6.765 2.05 ;
      POLYGON 6.205 1.32 5.765 1.32 5.765 0.48 5.325 0.48 5.325 0.36 5.885 0.36 5.885 1.2 6.205 1.2 ;
      POLYGON 5.725 1.64 5.485 1.64 5.485 1.52 5.525 1.52 5.525 1.28 4.115 1.28 4.115 1.11 3.095 1.11 3.095 1.14 2.855 1.14 2.855 1.02 2.975 1.02 2.975 0.99 4.235 0.99 4.235 1.16 5.525 1.16 5.525 0.62 5.645 0.62 5.645 1.52 5.725 1.52 ;
      POLYGON 5.225 0.86 5.135 0.86 5.135 1.04 4.355 1.04 4.355 0.8 4.235 0.8 4.235 0.68 4.475 0.68 4.475 0.92 5.015 0.92 5.015 0.74 5.105 0.74 5.105 0.62 5.225 0.62 ;
      RECT 3.555 1.64 5.125 1.76 ;
      POLYGON 4.895 0.8 4.655 0.8 4.655 0.56 4.115 0.56 4.115 0.72 3.795 0.72 3.795 0.8 3.555 0.8 3.555 0.68 3.675 0.68 3.675 0.6 3.995 0.6 3.995 0.44 4.775 0.44 4.775 0.68 4.895 0.68 ;
      POLYGON 3.875 0.48 3.555 0.48 3.555 0.56 2.775 0.56 2.775 0.86 2.735 0.86 2.735 1.57 2.775 1.57 2.775 1.81 2.655 1.81 2.655 1.69 2.615 1.69 2.615 0.74 2.655 0.74 2.655 0.56 2.555 0.56 2.555 0.53 2.145 0.53 2.145 1.13 1.805 1.13 1.805 1.2 1.565 1.2 1.565 1.01 2.025 1.01 2.025 0.41 2.675 0.41 2.675 0.44 3.435 0.44 3.435 0.36 3.875 0.36 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END SDFFSRX1

MACRO CLKAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X2 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.084 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 1.235 0.355 1.475 ;
        RECT 0.07 1.235 0.355 1.435 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.084 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.775 1.175 1.09 1.295 ;
        RECT 0.775 1.055 0.895 1.295 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 0.885 1.67 1.145 ;
        RECT 1.45 0.575 1.57 1.445 ;
        RECT 1.355 1.325 1.475 2.045 ;
        RECT 1.355 0.455 1.475 0.695 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 1.775 -0.18 1.895 0.695 ;
        RECT 0.875 -0.18 0.995 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 1.395 1.895 2.79 ;
        RECT 0.935 1.555 1.055 2.79 ;
        RECT 0.135 2.195 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.33 1.205 1.21 1.205 1.21 0.935 0.635 0.935 0.635 1.795 0.515 1.795 0.515 0.86 0.175 0.86 0.175 0.74 0.635 0.74 0.635 0.815 1.33 0.815 ;
  END
END CLKAND2X2

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.41 1.38 1.725 ;
        RECT 1.21 1.24 1.33 1.535 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 0.965 1.67 1.44 ;
        RECT 1.52 0.985 1.67 1.435 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.06 0.51 1.435 ;
        RECT 0.24 1.05 0.48 1.24 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.085 0.82 1.5 ;
        RECT 0.7 1.07 0.82 1.5 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3489 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 0.725 1.515 0.845 ;
        RECT 1.395 0.605 1.515 0.845 ;
        RECT 0.97 1 1.335 1.12 ;
        RECT 1.215 0.725 1.335 1.12 ;
        RECT 0.97 1 1.09 2.21 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 0.495 0.52 0.735 0.64 ;
        RECT 0.495 -0.18 0.615 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.71 1.56 1.83 2.79 ;
        RECT 0.22 1.56 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 0.7 1.815 0.7 1.815 0.485 1.095 0.485 1.095 0.88 0.135 0.88 0.135 0.64 0.255 0.64 0.255 0.76 0.975 0.76 0.975 0.365 1.935 0.365 ;
  END
END OAI22X1

MACRO OAI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.04 1.38 1.51 ;
        RECT 1.23 1.04 1.35 1.54 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.465 1.025 1.66 ;
        RECT 0.905 1.42 1.025 1.66 ;
        RECT 0.65 1.465 0.8 1.725 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.325 0.51 1.78 ;
        RECT 0.385 1.3 0.505 1.78 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 1.465 1.67 1.725 ;
        RECT 1.5 0.8 1.62 1.78 ;
        RECT 1.485 0.68 1.605 0.92 ;
        RECT 1.145 1.66 1.62 1.78 ;
        RECT 1.065 1.78 1.265 1.9 ;
        RECT 1.065 1.78 1.185 2.02 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.645 -0.18 0.765 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.485 1.9 1.605 2.79 ;
        RECT 0.425 1.9 0.545 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.185 0.92 1.11 0.92 1.11 1.16 0.225 1.16 0.225 0.68 0.345 0.68 0.345 1.04 0.99 1.04 0.99 0.8 1.065 0.8 1.065 0.68 1.185 0.68 ;
  END
END OAI21XL

MACRO DFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX2 0 0 ;
  SIZE 13.05 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 1.02 0.405 1.26 ;
        RECT 0.07 1.02 0.405 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.26 1.535 1.45 ;
        RECT 1.175 1.23 1.435 1.45 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8976 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.48 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.2 3.175 1.47 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.165 1.12 10.425 1.38 ;
        RECT 10.175 1.02 10.415 1.38 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.915 0.68 11.035 2.03 ;
        RECT 10.8 1.465 11.035 1.725 ;
        RECT 10.83 1.38 11.035 1.725 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.715 0.74 12.055 0.86 ;
        RECT 11.755 1.32 11.875 2.03 ;
        RECT 11.67 1.175 11.835 1.435 ;
        RECT 11.715 0.74 11.835 1.44 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.05 0.18 ;
        RECT 12.295 -0.18 12.535 0.32 ;
        RECT 11.335 -0.18 11.575 0.32 ;
        RECT 10.375 -0.18 10.615 0.32 ;
        RECT 9.265 -0.18 9.385 0.83 ;
        RECT 2.595 0.72 2.835 0.84 ;
        RECT 2.595 -0.18 2.715 0.84 ;
        RECT 1.435 -0.18 1.555 0.38 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.05 2.79 ;
        RECT 12.175 1.38 12.295 2.79 ;
        RECT 11.335 1.38 11.455 2.79 ;
        RECT 10.495 1.5 10.615 2.79 ;
        RECT 9.185 2.13 9.305 2.79 ;
        RECT 9.065 2.13 9.305 2.25 ;
        RECT 6.385 1.88 6.625 2 ;
        RECT 6.385 1.88 6.505 2.79 ;
        RECT 4.165 2 4.405 2.12 ;
        RECT 4.165 2 4.285 2.79 ;
        RECT 2.905 2.13 3.025 2.79 ;
        RECT 1.195 1.87 1.315 2.79 ;
        RECT 0.135 1.98 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.975 0.86 12.855 0.86 12.855 1.2 12.715 1.2 12.715 1.62 12.595 1.62 12.595 1.2 11.955 1.2 11.955 1.08 12.735 1.08 12.735 0.74 12.975 0.74 ;
      POLYGON 12.895 0.52 12.775 0.52 12.775 0.56 11.275 0.56 11.275 1.26 11.155 1.26 11.155 0.56 10.775 0.56 10.775 1.26 10.655 1.26 10.655 0.6 9.805 0.6 9.805 1.59 9.785 1.59 9.785 2.01 9.665 2.01 9.665 1.47 9.685 1.47 9.685 1.11 8.625 1.11 8.625 0.99 9.685 0.99 9.685 0.48 10.655 0.48 10.655 0.44 12.655 0.44 12.655 0.4 12.895 0.4 ;
      POLYGON 10.255 0.84 10.045 0.84 10.045 1.62 10.195 1.62 10.195 2.25 9.425 2.25 9.425 2.01 6.985 2.01 6.985 1.52 6.165 1.52 6.165 1.4 7.105 1.4 7.105 1.89 9.545 1.89 9.545 2.13 10.075 2.13 10.075 1.74 9.925 1.74 9.925 0.72 10.255 0.72 ;
      POLYGON 9.565 1.35 7.465 1.35 7.465 1.04 5.645 1.04 5.645 1.64 5.605 1.64 5.605 1.76 5.485 1.76 5.485 1.52 5.525 1.52 5.525 0.62 5.645 0.62 5.645 0.92 7.585 0.92 7.585 1.23 9.565 1.23 ;
      POLYGON 9.025 0.77 8.725 0.77 8.725 0.53 8.185 0.53 8.185 0.77 7.945 0.77 7.945 0.65 8.065 0.65 8.065 0.41 8.845 0.41 8.845 0.65 9.025 0.65 ;
      POLYGON 8.945 2.25 6.745 2.25 6.745 1.76 6.265 1.76 6.265 2 5.705 2 5.705 2.24 4.525 2.24 4.525 1.88 4.045 1.88 4.045 2.25 3.165 2.25 3.165 2.13 3.925 2.13 3.925 1.76 4.645 1.76 4.645 2.12 5.585 2.12 5.585 1.88 6.145 1.88 6.145 1.64 6.865 1.64 6.865 2.13 8.945 2.13 ;
      POLYGON 8.825 1.77 7.225 1.77 7.225 1.28 6.025 1.28 6.025 1.76 5.905 1.76 5.905 1.16 7.345 1.16 7.345 1.65 8.825 1.65 ;
      POLYGON 8.605 0.77 8.425 0.77 8.425 1.01 7.705 1.01 7.705 0.8 5.885 0.8 5.885 0.68 7.825 0.68 7.825 0.89 8.305 0.89 8.305 0.65 8.605 0.65 ;
      POLYGON 5.845 0.48 5.405 0.48 5.405 1.3 5.365 1.3 5.365 2 4.765 2 4.765 1.64 3.805 1.64 3.805 2.01 2.585 2.01 2.585 2.23 2.495 2.23 2.495 2.25 2.255 2.25 2.255 2.23 1.935 2.23 1.935 1.23 1.775 1.23 1.775 1.11 1.055 1.11 1.055 0.99 1.195 0.99 1.195 0.49 0.685 0.49 0.685 0.8 0.695 0.8 0.695 1.58 0.575 1.58 0.575 0.92 0.565 0.92 0.565 0.37 1.315 0.37 1.315 0.99 1.895 0.99 1.895 1.04 2.055 1.04 2.055 2.11 2.465 2.11 2.465 1.89 3.685 1.89 3.685 1.52 4.885 1.52 4.885 1.88 5.245 1.88 5.245 1.18 5.285 1.18 5.285 0.36 5.845 0.36 ;
      POLYGON 5.165 1.06 5.125 1.06 5.125 1.76 5.005 1.76 5.005 1.4 3.445 1.4 3.445 1.65 3.565 1.65 3.565 1.77 3.325 1.77 3.325 1.71 2.655 1.71 2.655 1.29 2.775 1.29 2.775 1.59 3.325 1.59 3.325 1.28 3.655 1.28 3.655 0.92 3.605 0.92 3.605 0.66 3.725 0.66 3.725 0.8 3.775 0.8 3.775 1.28 5.005 1.28 5.005 0.94 5.045 0.94 5.045 0.62 5.165 0.62 ;
      POLYGON 4.145 0.9 4.025 0.9 4.025 0.54 3.485 0.54 3.485 0.72 3.365 0.72 3.365 0.84 3.125 0.84 3.125 0.72 3.245 0.72 3.245 0.6 3.365 0.6 3.365 0.42 4.145 0.42 ;
      POLYGON 3.535 1.16 3.295 1.16 3.295 1.08 2.295 1.08 2.295 1.99 2.175 1.99 2.175 0.92 2.015 0.92 2.015 0.66 2.135 0.66 2.135 0.8 2.295 0.8 2.295 0.96 3.415 0.96 3.415 1.04 3.535 1.04 ;
      POLYGON 1.815 1.69 0.935 1.69 0.935 1.82 0.895 1.82 0.895 2.09 0.775 2.09 0.775 1.7 0.815 1.7 0.815 0.73 0.955 0.73 0.955 0.61 1.075 0.61 1.075 0.85 0.935 0.85 0.935 1.57 1.695 1.57 1.695 1.41 1.815 1.41 ;
  END
END DFFSRX2

MACRO OAI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.075 0.815 2.25 1.215 ;
        RECT 2.075 0.815 2.195 1.225 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 1.05 1.11 1.475 ;
        RECT 0.94 1.355 1.09 1.76 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.35 1.67 1.725 ;
        RECT 1.535 1.235 1.655 1.725 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.45 0.8 1.87 ;
        RECT 0.65 1.135 0.77 1.87 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.33 1.045 0.51 1.435 ;
        RECT 0.33 1.035 0.45 1.435 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4268 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.27 0.995 1.935 1.115 ;
        RECT 1.815 0.645 1.935 1.115 ;
        RECT 1.27 0.995 1.39 2.205 ;
        RECT 1.23 1.175 1.39 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 0.915 0.515 1.155 0.635 ;
        RECT 0.915 -0.18 1.035 0.635 ;
        RECT 0.135 -0.18 0.255 0.695 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 2.035 1.555 2.155 2.79 ;
        RECT 0.17 1.555 0.29 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.355 0.695 2.235 0.695 2.235 0.525 1.515 0.525 1.515 0.875 0.555 0.875 0.555 0.635 0.675 0.635 0.675 0.755 1.395 0.755 1.395 0.405 2.355 0.405 ;
  END
END OAI32X1

MACRO TLATNCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX6 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 1.14 0.565 1.52 ;
        RECT 0.305 1.165 0.565 1.38 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.465 1.145 1.67 ;
        RECT 0.935 1.36 1.055 1.71 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.285 1.34 7.405 2.12 ;
        RECT 7.265 0.405 7.385 1.04 ;
        RECT 7.105 1.34 7.405 1.46 ;
        RECT 7.085 0.92 7.385 1.04 ;
        RECT 7.105 0.92 7.225 1.46 ;
        RECT 5.605 1.04 7.225 1.16 ;
        RECT 6.445 1.04 6.565 2.12 ;
        RECT 6.425 0.405 6.545 1.16 ;
        RECT 5.525 0.885 5.73 1.04 ;
        RECT 5.605 0.885 5.725 2.12 ;
        RECT 5.525 0.4 5.645 1.04 ;
        RECT 5.58 1.04 7.225 1.145 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.845 -0.18 6.965 0.92 ;
        RECT 6.005 -0.18 6.125 0.92 ;
        RECT 5.105 -0.18 5.225 0.73 ;
        RECT 3.705 0.45 3.945 0.57 ;
        RECT 3.825 -0.18 3.945 0.57 ;
        RECT 2.245 -0.18 2.365 0.38 ;
        RECT 0.615 -0.18 0.735 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.865 1.34 6.985 2.79 ;
        RECT 6.025 1.34 6.145 2.79 ;
        RECT 5.185 1.77 5.305 2.79 ;
        RECT 4.345 1.77 4.465 2.79 ;
        RECT 3.445 2.23 3.565 2.79 ;
        RECT 2.055 2.25 2.295 2.79 ;
        RECT 0.755 1.83 0.875 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.405 1.24 5.305 1.24 5.305 1.65 4.885 1.65 4.885 2.08 4.765 2.08 4.765 1.65 4.045 1.65 4.045 2.08 3.925 2.08 3.925 1.53 5.185 1.53 5.185 0.97 4.545 0.97 4.545 0.81 4.465 0.81 4.465 0.57 4.585 0.57 4.585 0.69 4.665 0.69 4.665 0.85 5.405 0.85 ;
      POLYGON 5.065 1.41 3.765 1.41 3.765 1.05 3.225 1.05 3.225 1.37 3.105 1.37 3.105 1.87 2.985 1.87 2.985 1.37 2.055 1.37 2.055 1.25 3.105 1.25 3.105 0.65 3.345 0.65 3.345 0.77 3.225 0.77 3.225 0.93 3.885 0.93 3.885 1.29 4.945 1.29 4.945 1.09 5.065 1.09 ;
      POLYGON 4.425 1.17 4.305 1.17 4.305 1.05 4.225 1.05 4.225 0.81 3.465 0.81 3.465 0.53 2.985 0.53 2.985 0.78 2.845 0.78 2.845 1.13 1.935 1.13 1.935 1.73 2.645 1.73 2.645 1.77 2.775 1.77 2.775 1.89 2.525 1.89 2.525 1.85 1.815 1.85 1.815 1.25 1.755 1.25 1.755 1.01 2.725 1.01 2.725 0.66 2.865 0.66 2.865 0.41 3.585 0.41 3.585 0.69 4.345 0.69 4.345 0.93 4.425 0.93 ;
      POLYGON 3.585 1.29 3.465 1.29 3.465 2.11 3.2 2.11 3.2 2.13 2.285 2.13 2.285 2.09 1.415 2.09 1.415 1.85 1.275 1.85 1.275 0.66 1.395 0.66 1.395 1.73 1.535 1.73 1.535 1.97 2.405 1.97 2.405 2.01 3.08 2.01 3.08 1.99 3.345 1.99 3.345 1.17 3.585 1.17 ;
      POLYGON 2.745 0.5 2.605 0.5 2.605 0.62 2.005 0.62 2.005 0.54 1.635 0.54 1.635 1.37 1.695 1.37 1.695 1.61 1.575 1.61 1.575 1.49 1.515 1.49 1.515 0.54 1.155 0.54 1.155 1.24 1.035 1.24 1.035 1.02 0.185 1.02 0.185 1.64 0.455 1.64 0.455 1.95 0.335 1.95 0.335 1.76 0.065 1.76 0.065 0.78 0.135 0.78 0.135 0.66 0.255 0.66 0.255 0.9 1.035 0.9 1.035 0.42 2.125 0.42 2.125 0.5 2.485 0.5 2.485 0.38 2.745 0.38 ;
  END
END TLATNCAX6

MACRO OA22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 1.02 1.16 1.33 ;
        RECT 0.94 1.12 1.09 1.435 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.98 0.51 1.435 ;
        RECT 0.36 0.98 0.48 1.74 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.08 0.82 1.52 ;
        RECT 0.65 1.08 0.82 1.5 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.27 1.67 1.725 ;
        RECT 1.535 1.26 1.655 1.74 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.465 2.765 1.605 ;
        RECT 2.645 0.68 2.765 1.605 ;
        RECT 1.975 1.8 2.54 1.92 ;
        RECT 2.39 1.465 2.54 1.92 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 2.165 -0.18 2.285 0.4 ;
        RECT 0.615 -0.18 0.735 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.615 1.86 1.735 2.79 ;
        RECT 0.335 1.86 0.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.075 1.16 1.79 1.16 1.79 1.14 1.4 1.14 1.4 1.675 1.155 1.675 1.155 1.92 0.915 1.92 0.915 1.8 1.035 1.8 1.035 1.555 1.28 1.555 1.28 0.78 1.395 0.78 1.395 0.66 1.515 0.66 1.515 0.9 1.4 0.9 1.4 1.02 1.91 1.02 1.91 1.04 2.075 1.04 ;
      POLYGON 1.935 0.9 1.815 0.9 1.815 0.54 1.095 0.54 1.095 0.9 0.975 0.9 0.975 0.84 0.075 0.84 0.075 0.72 0.975 0.72 0.975 0.42 1.935 0.42 ;
  END
END OA22XL

MACRO AND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X8 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.65 0.94 1.77 1.235 ;
        RECT 0.595 0.94 1.77 1.06 ;
        RECT 0.63 0.94 0.87 1.175 ;
        RECT 0.595 0.94 0.87 1.09 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.18 1.435 1.45 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.95 1.295 5.07 2.21 ;
        RECT 4.81 0.715 5.05 0.835 ;
        RECT 2.43 1.295 5.07 1.415 ;
        RECT 2.35 0.765 4.93 0.885 ;
        RECT 4.13 0.765 4.28 1.145 ;
        RECT 4.13 0.715 4.25 1.415 ;
        RECT 4.11 1.295 4.23 2.21 ;
        RECT 3.97 0.715 4.25 0.885 ;
        RECT 3.27 1.295 3.39 2.21 ;
        RECT 3.13 0.715 3.37 0.885 ;
        RECT 2.43 1.295 2.55 2.21 ;
        RECT 2.23 0.715 2.47 0.835 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 4.45 -0.18 4.57 0.645 ;
        RECT 3.61 -0.18 3.73 0.645 ;
        RECT 2.71 -0.18 2.83 0.64 ;
        RECT 1.81 0.46 2.05 0.58 ;
        RECT 1.81 -0.18 1.93 0.58 ;
        RECT 0.53 -0.18 0.65 0.705 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.53 1.535 4.65 2.79 ;
        RECT 3.69 1.535 3.81 2.79 ;
        RECT 2.85 1.535 2.97 2.79 ;
        RECT 2.01 1.81 2.13 2.79 ;
        RECT 1.17 1.81 1.29 2.79 ;
        RECT 0.33 1.56 0.45 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.01 1.175 2.01 1.175 2.01 1.69 1.71 1.69 1.71 2.21 1.59 2.21 1.59 1.69 0.87 1.69 0.87 2.21 0.75 2.21 0.75 1.56 0.87 1.56 0.87 1.57 1.59 1.57 1.59 1.56 1.71 1.56 1.71 1.57 1.89 1.57 1.89 0.82 1.11 0.82 1.11 0.7 2.01 0.7 2.01 1.055 4.01 1.055 ;
  END
END AND2X8

MACRO TLATNX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX4 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.93 0.855 1.14 ;
        RECT 0.555 1.02 0.795 1.2 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.77 1.345 8.92 1.76 ;
        RECT 8.795 1.12 8.915 1.76 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.295 1.32 2.415 2.21 ;
        RECT 1.52 1.32 2.415 1.44 ;
        RECT 1.095 0.8 2.175 0.92 ;
        RECT 2.055 0.68 2.175 0.92 ;
        RECT 1.55 0.8 1.67 1.56 ;
        RECT 1.455 1.44 1.575 2.21 ;
        RECT 1.52 1.175 1.67 1.56 ;
        RECT 1.095 0.68 1.215 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.935 0.8 6.015 0.92 ;
        RECT 5.895 0.68 6.015 0.92 ;
        RECT 5.655 1.52 5.775 2.21 ;
        RECT 4.945 1.52 5.775 1.64 ;
        RECT 4.815 1.55 5.205 1.67 ;
        RECT 5.085 0.8 5.205 1.67 ;
        RECT 4.935 0.68 5.055 0.92 ;
        RECT 4.815 1.55 4.935 2.21 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.735 -0.18 8.855 0.4 ;
        RECT 7.335 -0.18 7.455 0.4 ;
        RECT 6.315 -0.18 6.555 0.32 ;
        RECT 5.355 -0.18 5.595 0.32 ;
        RECT 4.395 -0.18 4.635 0.32 ;
        RECT 3.435 -0.18 3.675 0.32 ;
        RECT 2.475 -0.18 2.715 0.32 ;
        RECT 1.515 -0.18 1.755 0.32 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.755 1.88 8.875 2.79 ;
        RECT 6.915 1.66 7.155 2.06 ;
        RECT 6.915 1.66 7.035 2.79 ;
        RECT 6.075 1.56 6.195 2.79 ;
        RECT 5.235 1.79 5.355 2.79 ;
        RECT 4.395 1.56 4.515 2.79 ;
        RECT 3.555 1.56 3.675 2.79 ;
        RECT 2.715 1.56 2.835 2.79 ;
        RECT 1.875 1.56 1.995 2.79 ;
        RECT 1.035 1.56 1.155 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.455 0.86 9.335 0.86 9.335 1 9.295 1 9.295 2 9.175 2 9.175 1 8.635 1 8.635 1.4 8.395 1.4 8.395 0.88 9.215 0.88 9.215 0.74 9.455 0.74 ;
      POLYGON 9.235 0.52 9.095 0.52 9.095 0.64 8.495 0.64 8.495 0.62 7.855 0.62 7.855 1.5 7.975 1.5 7.975 1.62 7.735 1.62 7.735 0.64 7.095 0.64 7.095 0.56 0.975 0.56 0.975 0.68 0.255 0.68 0.255 1.32 0.575 1.32 0.575 1.8 0.455 1.8 0.455 1.44 0.135 1.44 0.135 0.56 0.855 0.56 0.855 0.44 7.215 0.44 7.215 0.52 7.735 0.52 7.735 0.5 8.135 0.5 8.135 0.4 8.375 0.4 8.375 0.5 8.615 0.5 8.615 0.52 8.975 0.52 8.975 0.4 9.235 0.4 ;
      POLYGON 8.215 2 8.095 2 8.095 1.86 7.495 1.86 7.495 1.5 6.815 1.5 6.815 1.26 6.935 1.26 6.935 1.38 7.615 1.38 7.615 1.74 8.095 1.74 8.095 0.86 7.975 0.86 7.975 0.74 8.215 0.74 ;
      POLYGON 7.555 1.26 7.435 1.26 7.435 1.14 6.675 1.14 6.675 2.12 6.555 2.12 6.555 1.26 5.695 1.26 5.695 1.14 6.555 1.14 6.555 1.02 6.855 1.02 6.855 0.68 6.975 0.68 6.975 1.02 7.555 1.02 ;
      POLYGON 4.095 0.92 3.255 0.92 3.255 1.32 4.095 1.32 4.095 2.21 3.975 2.21 3.975 1.44 3.255 1.44 3.255 2.21 3.135 2.21 3.135 1.2 2.095 1.2 2.095 1.08 3.135 1.08 3.135 0.92 3.015 0.92 3.015 0.68 3.135 0.68 3.135 0.8 3.975 0.8 3.975 0.68 4.095 0.68 ;
  END
END TLATNX4

MACRO SMDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX8 0 0 ;
  SIZE 14.21 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.445 2.775 2.19 ;
        RECT 2.655 0.665 2.775 0.905 ;
        RECT 2.635 0.785 2.755 1.565 ;
        RECT 0.07 0.905 2.755 1.025 ;
        RECT 1.815 0.665 1.935 2.19 ;
        RECT 0.975 0.665 1.095 2.185 ;
        RECT 0.135 0.665 0.255 2.185 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 1.175 5.205 1.38 ;
        RECT 5.085 1.03 5.205 1.38 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.67 1.16 9.915 1.28 ;
        RECT 9.67 0.885 9.79 1.28 ;
        RECT 9.64 0.885 9.79 1.145 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.38 0.885 11.53 1.145 ;
        RECT 11.295 1.025 11.415 1.385 ;
    END
  END SE
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.595 1.265 11.835 1.385 ;
        RECT 11.67 0.885 11.82 1.145 ;
        RECT 11.67 0.885 11.79 1.385 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.05 1.21 13.355 1.42 ;
        RECT 13.05 1.21 13.325 1.445 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.495 0.97 13.615 1.21 ;
        RECT 12.535 0.97 13.615 1.09 ;
        RECT 12.775 0.94 13.035 1.09 ;
        RECT 12.315 1 12.655 1.12 ;
        RECT 12.195 1.265 12.435 1.385 ;
        RECT 12.315 1 12.435 1.385 ;
    END
  END S0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.21 0.18 ;
        RECT 13.335 -0.18 13.455 0.82 ;
        RECT 12.055 -0.18 12.175 0.64 ;
        RECT 9.855 -0.18 9.975 0.765 ;
        RECT 7.585 0.41 7.825 0.53 ;
        RECT 7.705 -0.18 7.825 0.53 ;
        RECT 5.325 0.31 5.565 0.43 ;
        RECT 5.445 -0.18 5.565 0.43 ;
        RECT 3.915 -0.18 4.035 0.65 ;
        RECT 3.075 -0.18 3.195 0.65 ;
        RECT 2.235 -0.18 2.355 0.655 ;
        RECT 1.395 -0.18 1.515 0.655 ;
        RECT 0.555 -0.18 0.675 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.21 2.79 ;
        RECT 13.135 1.805 13.255 2.79 ;
        RECT 11.755 1.745 11.875 2.79 ;
        RECT 9.795 1.75 9.915 2.79 ;
        RECT 7.585 2.01 7.825 2.13 ;
        RECT 7.585 2.01 7.705 2.79 ;
        RECT 5.685 1.98 5.805 2.79 ;
        RECT 3.915 1.54 4.035 2.79 ;
        RECT 3.075 1.54 3.195 2.79 ;
        RECT 2.235 1.445 2.355 2.79 ;
        RECT 1.395 1.445 1.515 2.79 ;
        RECT 0.555 1.445 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.875 0.82 13.855 0.82 13.855 1.685 13.775 1.685 13.775 1.805 13.655 1.805 13.655 1.685 12.635 1.685 12.635 1.24 12.755 1.24 12.755 1.565 13.735 1.565 13.735 0.7 13.755 0.7 13.755 0.58 13.875 0.58 ;
      POLYGON 12.815 0.82 12.415 0.82 12.415 0.88 12.075 0.88 12.075 1.505 12.515 1.505 12.515 2.21 12.395 2.21 12.395 1.625 11.035 1.625 11.035 1.82 10.915 1.82 10.915 1.49 11.055 1.49 11.055 0.765 11.035 0.765 11.035 0.645 11.275 0.645 11.275 0.765 11.175 0.765 11.175 1.505 11.955 1.505 11.955 0.76 12.295 0.76 12.295 0.7 12.695 0.7 12.695 0.56 12.815 0.56 ;
      POLYGON 11.715 0.765 11.475 0.765 11.475 0.525 10.915 0.525 10.915 0.885 10.935 0.885 10.935 1.37 10.795 1.37 10.795 1.97 11.395 1.97 11.395 2.21 11.275 2.21 11.275 2.09 10.675 2.09 10.675 1.27 10.395 1.27 10.395 1.39 10.275 1.39 10.275 1.15 10.815 1.15 10.815 1.005 10.795 1.005 10.795 0.405 11.595 0.405 11.595 0.645 11.715 0.645 ;
      POLYGON 10.675 0.77 10.555 0.77 10.555 1.005 10.155 1.005 10.155 1.51 10.555 1.51 10.555 2.14 10.435 2.14 10.435 1.63 9.105 1.63 9.105 1.93 8.985 1.93 8.985 1.44 9.025 1.44 9.025 0.72 8.985 0.72 8.985 0.6 9.225 0.6 9.225 0.72 9.145 0.72 9.145 1.51 10.035 1.51 10.035 0.885 10.435 0.885 10.435 0.65 10.675 0.65 ;
      POLYGON 9.555 0.765 9.435 0.765 9.435 0.48 8.865 0.48 8.865 1.08 8.905 1.08 8.905 1.32 8.865 1.32 8.865 2.05 9.315 2.05 9.315 1.93 9.555 1.93 9.555 2.05 9.435 2.05 9.435 2.17 8.745 2.17 8.745 0.48 8.265 0.48 8.265 0.92 8.385 0.92 8.385 1.04 8.145 1.04 8.145 0.77 7.345 0.77 7.345 0.48 6.865 0.48 6.865 0.84 6.985 0.84 6.985 1.12 6.865 1.12 6.865 0.96 6.745 0.96 6.745 0.36 7.465 0.36 7.465 0.65 8.145 0.65 8.145 0.36 9.555 0.36 ;
      POLYGON 8.625 1.93 8.505 1.93 8.505 1.28 7.485 1.28 7.485 1.25 7.365 1.25 7.365 1.13 7.605 1.13 7.605 1.16 8.505 1.16 8.505 0.72 8.385 0.72 8.385 0.6 8.625 0.6 ;
      POLYGON 8.345 2.25 8.225 2.25 8.225 1.89 7.285 1.89 7.285 2.17 5.945 2.17 5.945 0.91 4.825 0.91 4.825 1.5 5.305 1.5 5.305 1.62 4.705 1.62 4.705 0.6 4.965 0.6 4.965 0.79 6.065 0.79 6.065 2.05 6.625 2.05 6.625 1.32 6.525 1.32 6.525 1.08 6.645 1.08 6.645 1.2 6.745 1.2 6.745 2.05 7.165 2.05 7.165 1.77 8.345 1.77 ;
      POLYGON 8.025 1.04 7.725 1.04 7.725 1.01 7.225 1.01 7.225 1.65 7.105 1.65 7.105 0.72 6.985 0.72 6.985 0.6 7.225 0.6 7.225 0.89 7.845 0.89 7.845 0.92 8.025 0.92 ;
      POLYGON 6.505 1.93 6.385 1.93 6.385 1.56 6.285 1.56 6.285 0.67 5.085 0.67 5.085 0.48 4.275 0.48 4.275 1.18 4.155 1.18 4.155 0.36 5.205 0.36 5.205 0.55 6.285 0.55 6.285 0.54 6.405 0.54 6.405 1.44 6.505 1.44 ;
      POLYGON 5.725 1.86 4.455 1.86 4.455 2.19 4.335 2.19 4.335 1.54 4.395 1.54 4.395 1.42 3.615 1.42 3.615 2.19 3.495 2.19 3.495 1.225 2.875 1.225 2.875 1.105 3.495 1.105 3.495 0.6 3.615 0.6 3.615 1.3 4.395 1.3 4.395 0.6 4.515 0.6 4.515 1.74 5.605 1.74 5.605 1.07 5.725 1.07 ;
  END
END SMDFFHQX8

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.97 1.055 1.21 1.195 ;
        RECT 0.94 1.15 1.09 1.435 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.02 0.82 1.435 ;
        RECT 0.7 1.005 0.82 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.825 0.51 1.28 ;
        RECT 0.38 0.825 0.5 1.305 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3196 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 0.885 1.67 1.145 ;
        RECT 1.395 0.765 1.515 2.21 ;
        RECT 0.86 0.765 1.515 0.885 ;
        RECT 0.86 0.645 0.98 0.885 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 1.22 0.525 1.46 0.645 ;
        RECT 1.22 -0.18 1.34 0.645 ;
        RECT 0.22 -0.18 0.34 0.705 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.555 1.795 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.095 2.21 0.975 2.21 0.975 1.675 0.255 1.675 0.255 2.21 0.135 2.21 0.135 1.555 1.095 1.555 ;
  END
END AOI21X1

MACRO DFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX4 0 0 ;
  SIZE 10.73 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.165 1.1 0.355 1.34 ;
        RECT 0.07 1.175 0.285 1.435 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 1.1 0.8 1.525 ;
        RECT 0.665 1.08 0.795 1.525 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.185 1.725 1.38 ;
        RECT 1.465 1.02 1.585 1.38 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.575 0.74 7.775 0.86 ;
        RECT 7.635 1.44 7.755 2.21 ;
        RECT 7.455 1.44 7.755 1.56 ;
        RECT 6.77 1.32 7.575 1.44 ;
        RECT 6.795 0.74 6.915 2.21 ;
        RECT 6.74 1.175 6.915 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.495 0.74 9.695 0.86 ;
        RECT 9.315 1.32 9.435 2.21 ;
        RECT 8.48 1.32 9.435 1.44 ;
        RECT 8.51 0.74 8.63 1.56 ;
        RECT 8.475 1.44 8.595 2.21 ;
        RECT 8.48 1.175 8.63 1.56 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.73 0.18 ;
        RECT 10.055 -0.18 10.175 0.73 ;
        RECT 8.975 -0.18 9.215 0.38 ;
        RECT 8.015 -0.18 8.255 0.38 ;
        RECT 7.055 -0.18 7.295 0.38 ;
        RECT 6.095 -0.18 6.335 0.38 ;
        RECT 5.255 -0.18 5.375 0.92 ;
        RECT 3.605 -0.18 3.845 0.32 ;
        RECT 1.615 -0.18 1.735 0.66 ;
        RECT 0.165 -0.18 0.285 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.73 2.79 ;
        RECT 9.735 1.6 9.855 2.79 ;
        RECT 8.895 1.56 9.015 2.79 ;
        RECT 8.055 1.56 8.175 2.79 ;
        RECT 7.215 1.56 7.335 2.79 ;
        RECT 6.375 1.56 6.495 2.79 ;
        RECT 5.475 1.64 5.595 2.79 ;
        RECT 3.605 1.75 3.725 2.79 ;
        RECT 1.765 1.98 1.885 2.79 ;
        RECT 0.975 1.98 1.095 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.595 0.92 10.415 0.92 10.415 1.48 10.275 1.48 10.275 2.21 10.155 2.21 10.155 1.48 9.555 1.48 9.555 1.3 9.795 1.3 9.795 1.36 10.295 1.36 10.295 0.8 10.475 0.8 10.475 0.68 10.595 0.68 ;
      POLYGON 10.135 1.24 10.015 1.24 10.015 0.97 9.815 0.97 9.815 0.62 6.325 0.62 6.325 0.68 5.795 0.68 5.795 0.8 6.155 0.8 6.155 1.3 6.62 1.3 6.62 1.42 6.015 1.42 6.015 2.15 5.895 2.15 5.895 1.42 5.515 1.42 5.515 1.52 5.395 1.52 5.395 1.28 5.515 1.28 5.515 1.3 6.035 1.3 6.035 0.92 5.675 0.92 5.675 0.56 6.205 0.56 6.205 0.5 9.935 0.5 9.935 0.85 10.135 0.85 ;
      POLYGON 5.915 1.18 5.675 1.18 5.675 1.16 5.275 1.16 5.275 1.77 4.935 1.77 4.935 1.81 4.695 1.81 4.695 1.69 4.815 1.69 4.815 1.65 5.155 1.65 5.155 1.16 4.615 1.16 4.615 0.68 4.735 0.68 4.735 1.04 5.915 1.04 ;
      POLYGON 5.035 1.53 4.915 1.53 4.915 1.4 4.375 1.4 4.375 0.56 2.785 0.56 2.785 1.37 2.845 1.37 2.845 1.49 2.605 1.49 2.605 1.37 2.665 1.37 2.665 0.56 2.245 0.56 2.245 1.58 2.125 1.58 2.125 0.66 2.035 0.66 2.035 0.42 2.155 0.42 2.155 0.44 3.065 0.44 3.065 0.4 3.305 0.4 3.305 0.44 4.495 0.44 4.495 1.28 5.035 1.28 ;
      POLYGON 4.255 1.87 4.135 1.87 4.135 1.49 3.405 1.49 3.405 1.37 4.135 1.37 4.135 0.68 4.255 0.68 ;
      POLYGON 4.015 1.25 3.085 1.25 3.085 1.87 2.965 1.87 2.965 0.86 2.905 0.86 2.905 0.74 3.145 0.74 3.145 0.86 3.085 0.86 3.085 1.13 4.015 1.13 ;
      POLYGON 2.645 1.87 2.525 1.87 2.525 1.86 0.92 1.86 0.92 1.77 0.435 1.77 0.435 1.65 0.92 1.65 0.92 0.96 0.805 0.96 0.805 0.68 0.925 0.68 0.925 0.84 1.04 0.84 1.04 1.74 2.365 1.74 2.365 0.8 2.425 0.8 2.425 0.68 2.545 0.68 2.545 0.92 2.485 0.92 2.485 1.63 2.645 1.63 ;
      POLYGON 1.985 1.16 1.865 1.16 1.865 0.9 1.345 0.9 1.345 1.5 1.465 1.5 1.465 1.62 1.225 1.62 1.225 0.66 1.195 0.66 1.195 0.42 1.315 0.42 1.315 0.54 1.345 0.54 1.345 0.78 1.985 0.78 ;
  END
END DFFTRX4

MACRO TLATNCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX3 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 1.02 0.395 1.28 ;
        RECT 0.07 1.02 0.395 1.16 ;
        RECT 0.07 0.885 0.22 1.16 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.325 1.23 1.445 1.58 ;
        RECT 1.175 1.23 1.445 1.435 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.825 1.32 5.945 2.21 ;
        RECT 5.825 0.6 5.945 0.84 ;
        RECT 5 1.32 5.945 1.44 ;
        RECT 5.645 0.72 5.945 0.84 ;
        RECT 5 0.84 5.765 0.96 ;
        RECT 5 1.175 5.15 1.44 ;
        RECT 5 0.72 5.12 1.56 ;
        RECT 4.985 1.44 5.105 2.21 ;
        RECT 4.985 0.6 5.105 0.84 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.405 -0.18 5.525 0.65 ;
        RECT 4.505 0.47 4.745 0.59 ;
        RECT 4.505 -0.18 4.625 0.59 ;
        RECT 2.905 -0.18 3.025 0.38 ;
        RECT 1.425 -0.18 1.545 0.63 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.405 1.56 5.525 2.79 ;
        RECT 4.565 1.76 4.685 2.79 ;
        RECT 3.665 1.62 3.905 2.15 ;
        RECT 3.665 1.62 3.785 2.79 ;
        RECT 2.545 1.97 2.665 2.79 ;
        RECT 1.265 1.97 1.385 2.79 ;
        RECT 0.135 1.46 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.825 1.4 4.665 1.4 4.665 1.64 4.265 1.64 4.265 2.21 4.145 2.21 4.145 1.52 4.545 1.52 4.545 0.83 4.045 0.83 4.045 0.78 3.865 0.78 3.865 0.66 4.165 0.66 4.165 0.71 4.665 0.71 4.665 1.16 4.825 1.16 ;
      POLYGON 4.425 1.4 3.085 1.4 3.085 2.09 2.965 2.09 2.965 1.4 2.425 1.4 2.425 1.28 3.385 1.28 3.385 0.66 3.505 0.66 3.505 1.28 4.305 1.28 4.305 1.16 4.425 1.16 ;
      POLYGON 4.045 1.1 3.805 1.1 3.805 1.02 3.625 1.02 3.625 0.54 3.265 0.54 3.265 0.62 2.665 0.62 2.665 0.6 2.025 0.6 2.025 1.71 1.785 1.71 1.785 1.82 1.145 1.82 1.145 1.94 0.965 1.94 0.965 2.09 0.845 2.09 0.845 1.82 1.025 1.82 1.025 1.7 1.665 1.7 1.665 1.59 1.905 1.59 1.905 0.87 1.11 0.87 1.11 0.84 0.885 0.84 0.885 0.72 1.23 0.72 1.23 0.75 1.905 0.75 1.905 0.48 2.305 0.48 2.305 0.38 2.545 0.38 2.545 0.48 2.785 0.48 2.785 0.5 3.145 0.5 3.145 0.42 3.745 0.42 3.745 0.9 3.925 0.9 3.925 0.98 4.045 0.98 ;
      POLYGON 3.105 1.16 2.305 1.16 2.305 1.95 2.025 1.95 2.025 2.09 1.905 2.09 1.905 1.83 2.185 1.83 2.185 0.84 2.145 0.84 2.145 0.72 2.385 0.72 2.385 0.84 2.305 0.84 2.305 1.04 3.105 1.04 ;
      POLYGON 1.785 1.45 1.665 1.45 1.665 1.11 1.055 1.11 1.055 1.18 0.815 1.18 0.815 1.11 0.675 1.11 0.675 1.58 0.555 1.58 0.555 0.68 0.675 0.68 0.675 0.99 1.785 0.99 ;
  END
END TLATNCAX3

MACRO FILL4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL4 0 0 ;
  SIZE 1.16 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.16 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.16 0.18 ;
    END
  END VSS
END FILL4

MACRO OAI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.125 1.38 1.615 ;
        RECT 1.23 1.125 1.38 1.585 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.885 1.7 1.27 ;
        RECT 1.58 0.875 1.7 1.27 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.885 0.51 1.34 ;
        RECT 0.36 0.885 0.48 1.365 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.335 1.09 1.725 ;
        RECT 0.94 1.145 1.06 1.725 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 1.465 1.96 1.725 ;
        RECT 1.84 0.525 1.96 1.725 ;
        RECT 1.42 1.735 1.72 1.855 ;
        RECT 1.6 1.465 1.72 1.855 ;
        RECT 1.42 1.735 1.54 1.975 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1 -0.18 1.12 0.765 ;
        RECT 0.16 -0.18 0.28 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.84 1.845 1.96 2.79 ;
        RECT 0.46 1.845 0.58 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.6 0.705 1.4 0.705 1.4 1.005 0.63 1.005 0.63 0.765 0.58 0.765 0.58 0.525 0.7 0.525 0.7 0.645 0.75 0.645 0.75 0.885 1.28 0.885 1.28 0.585 1.6 0.585 ;
  END
END OAI31XL

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 1.45 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1 0.82 1.38 ;
        RECT 0.65 1.175 0.8 1.55 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.785 0.51 1.235 ;
        RECT 0.36 0.76 0.48 1.235 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3196 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.94 0.76 1.06 2.005 ;
        RECT 0.63 0.76 1.06 0.88 ;
        RECT 0.63 0.545 0.75 0.88 ;
        RECT 0.62 0.425 0.74 0.665 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.45 0.18 ;
        RECT 1.04 -0.18 1.16 0.64 ;
        RECT 0.2 -0.18 0.32 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.45 2.79 ;
        RECT 0.2 1.355 0.32 2.79 ;
    END
  END VDD
END NOR2X1

MACRO SDFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX4 0 0 ;
  SIZE 16.53 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.655 1.46 1.895 1.58 ;
        RECT 1.655 0.36 1.775 1.58 ;
        RECT 0.955 0.36 1.775 0.48 ;
        RECT 0.355 0.92 1.295 1.04 ;
        RECT 0.885 0.92 1.145 1.09 ;
        RECT 0.955 0.36 1.075 1.09 ;
        RECT 0.355 0.92 0.475 1.16 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.235 0.955 1.435 ;
        RECT 0.595 1.21 0.855 1.435 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 1.935 1.175 2.25 1.295 ;
        RECT 1.935 1.055 2.055 1.295 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.9 2.885 1.12 ;
        RECT 2.655 0.9 2.775 1.29 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.975 1.165 7.235 1.38 ;
        RECT 7.105 1 7.225 1.38 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 1.185 7.815 1.38 ;
        RECT 7.565 1 7.685 1.38 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.165 0.7 13.365 0.82 ;
        RECT 13.185 1.44 13.305 2.21 ;
        RECT 12.905 1.44 13.305 1.56 ;
        RECT 12.25 1.32 13.025 1.44 ;
        RECT 12.28 0.7 12.4 1.56 ;
        RECT 12.245 1.44 12.365 2.21 ;
        RECT 12.25 1.175 12.4 1.56 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.085 0.7 15.285 0.82 ;
        RECT 14.905 1.56 15.025 2.21 ;
        RECT 14.885 1.32 15.005 1.68 ;
        RECT 14.245 1.32 15.005 1.44 ;
        RECT 14.245 1.175 14.43 1.44 ;
        RECT 14.065 1.44 14.365 1.56 ;
        RECT 14.245 0.7 14.365 1.56 ;
        RECT 14.065 1.44 14.185 2.21 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 16.53 0.18 ;
        RECT 15.645 0.51 15.885 0.63 ;
        RECT 15.765 -0.18 15.885 0.63 ;
        RECT 14.565 -0.18 14.805 0.34 ;
        RECT 13.605 -0.18 13.845 0.34 ;
        RECT 12.645 -0.18 12.885 0.34 ;
        RECT 11.565 0.6 11.805 0.72 ;
        RECT 11.565 -0.18 11.685 0.72 ;
        RECT 10.785 -0.18 10.905 0.86 ;
        RECT 7.305 0.52 7.545 0.64 ;
        RECT 7.305 -0.18 7.425 0.64 ;
        RECT 4.705 -0.18 4.945 0.34 ;
        RECT 1.895 -0.18 2.015 0.78 ;
        RECT 0.615 -0.18 0.735 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 16.53 2.79 ;
        RECT 15.325 1.56 15.445 2.79 ;
        RECT 14.485 1.56 14.605 2.79 ;
        RECT 13.645 1.56 13.765 2.79 ;
        RECT 12.665 1.56 12.785 2.79 ;
        RECT 11.825 1.6 11.945 2.79 ;
        RECT 10.985 1.76 11.105 2.79 ;
        RECT 9.925 1.88 10.045 2.79 ;
        RECT 7.215 1.98 7.335 2.79 ;
        RECT 7.095 1.98 7.335 2.1 ;
        RECT 5.435 2.24 5.675 2.79 ;
        RECT 4.565 2.24 4.805 2.79 ;
        RECT 2.155 1.94 2.395 2.06 ;
        RECT 2.155 1.94 2.275 2.79 ;
        RECT 0.675 1.88 0.795 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 16.245 1.44 15.865 1.44 15.865 2.21 15.745 2.21 15.745 1.44 15.125 1.44 15.125 1.3 15.365 1.3 15.365 1.32 16.125 1.32 16.125 0.64 16.245 0.64 ;
      POLYGON 15.725 1.2 15.605 1.2 15.605 0.87 15.405 0.87 15.405 0.58 12.045 0.58 12.045 0.96 11.505 0.96 11.505 1.22 12.125 1.22 12.125 1.34 11.525 1.34 11.525 2.12 11.405 2.12 11.405 1.34 11.385 1.34 11.385 1.14 10.245 1.14 10.245 1.02 11.205 1.02 11.205 0.64 11.325 0.64 11.325 0.84 11.925 0.84 11.925 0.46 15.525 0.46 15.525 0.75 15.725 0.75 ;
      POLYGON 11.265 1.52 8.845 1.52 8.845 1.89 8.725 1.89 8.725 1.4 8.655 1.4 8.655 0.68 8.775 0.68 8.775 1.28 8.845 1.28 8.845 1.4 11.145 1.4 11.145 1.26 11.265 1.26 ;
      POLYGON 10.745 1.94 10.265 1.94 10.265 1.76 9.59 1.76 9.59 1.81 9.085 1.81 9.085 1.69 9.47 1.69 9.47 1.64 10.385 1.64 10.385 1.82 10.745 1.82 ;
      POLYGON 10.485 0.86 10.365 0.86 10.365 0.74 10.185 0.74 10.185 0.5 9.775 0.5 9.775 0.8 9.465 0.8 9.465 0.68 9.655 0.68 9.655 0.38 10.305 0.38 10.305 0.62 10.485 0.62 ;
      POLYGON 10.065 1.04 9.225 1.04 9.225 0.92 9.135 0.92 9.135 0.68 9.255 0.68 9.255 0.8 9.345 0.8 9.345 0.92 9.945 0.92 9.945 0.62 10.065 0.62 ;
      POLYGON 9.865 1.28 8.985 1.28 8.985 1.16 8.895 1.16 8.895 0.56 7.965 0.56 7.965 0.74 8.055 0.74 8.055 1.62 7.935 1.62 7.935 0.86 7.785 0.86 7.785 0.88 7.065 0.88 7.065 0.5 6.65 0.5 6.65 0.48 6.265 0.48 6.265 0.36 6.77 0.36 6.77 0.38 7.185 0.38 7.185 0.76 7.665 0.76 7.665 0.62 7.845 0.62 7.845 0.44 9.015 0.44 9.015 1.04 9.105 1.04 9.105 1.16 9.865 1.16 ;
      POLYGON 9.105 2.25 7.955 2.25 7.955 2.13 7.455 2.13 7.455 1.86 6.375 1.86 6.375 1.64 5.045 1.64 5.045 1.52 5.185 1.52 5.185 1 4.345 1 4.345 1.28 4.225 1.28 4.225 0.88 5.185 0.88 5.185 0.7 5.425 0.7 5.425 0.82 5.305 0.82 5.305 1.52 6.495 1.52 6.495 1.74 7.575 1.74 7.575 2.01 8.075 2.01 8.075 2.13 8.485 2.13 8.485 1.64 8.415 1.64 8.415 1.04 8.535 1.04 8.535 1.52 8.605 1.52 8.605 2.13 9.105 2.13 ;
      POLYGON 8.365 2.01 8.245 2.01 8.245 1.89 7.695 1.89 7.695 1.62 6.615 1.62 6.615 1.4 5.545 1.4 5.545 0.58 4.465 0.58 4.465 0.5 4.345 0.5 4.345 0.38 4.585 0.38 4.585 0.46 5.525 0.46 5.525 0.38 6.145 0.38 6.145 0.6 6.465 0.6 6.465 0.68 6.585 0.68 6.585 0.8 6.345 0.8 6.345 0.72 6.025 0.72 6.025 0.5 5.665 0.5 5.665 1.28 6.855 1.28 6.855 1.5 7.815 1.5 7.815 1.77 8.175 1.77 8.175 0.8 8.235 0.8 8.235 0.68 8.355 0.68 8.355 0.92 8.295 0.92 8.295 1.77 8.365 1.77 ;
      POLYGON 6.975 2.25 6.4 2.25 6.4 2.1 6.135 2.1 6.135 1.88 4.805 1.88 4.805 1.52 4.245 1.52 4.245 1.56 4.005 1.56 4.005 1.52 3.985 1.52 3.985 0.52 3.5 0.52 3.5 0.54 2.555 0.54 2.555 0.66 3.125 0.66 3.125 1.94 2.755 1.94 2.755 1.82 3.005 1.82 3.005 0.78 2.435 0.78 2.435 0.42 3.38 0.42 3.38 0.4 3.525 0.4 3.525 0.36 3.765 0.36 3.765 0.4 4.105 0.4 4.105 1.4 4.805 1.4 4.805 1.12 4.965 1.12 4.965 1.36 4.925 1.36 4.925 1.76 6.255 1.76 6.255 1.98 6.52 1.98 6.52 2.13 6.975 2.13 ;
      POLYGON 6.945 1.04 5.785 1.04 5.785 0.62 5.905 0.62 5.905 0.92 6.825 0.92 6.825 0.62 6.945 0.62 ;
      POLYGON 6.015 2.12 4.45 2.12 4.45 2.06 3.925 2.06 3.925 1.82 3.745 1.82 3.745 0.64 3.865 0.64 3.865 1.7 4.045 1.7 4.045 1.94 4.57 1.94 4.57 2 6.015 2 ;
      POLYGON 3.625 2.18 2.515 2.18 2.515 1.82 1.575 1.82 1.575 2 1.455 2 1.455 1.88 1.415 1.88 1.415 0.72 1.195 0.72 1.195 0.6 1.535 0.6 1.535 1.7 2.635 1.7 2.635 2.06 3.505 2.06 3.505 0.82 3.265 0.82 3.265 0.7 3.625 0.7 ;
      POLYGON 1.295 1.675 0.375 1.675 0.375 2 0.255 2 0.255 1.795 0.115 1.795 0.115 0.68 0.195 0.68 0.195 0.54 0.315 0.54 0.315 0.8 0.235 0.8 0.235 1.555 1.175 1.555 1.175 1.21 1.295 1.21 ;
  END
END SDFFSRX4

MACRO SMDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX2 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.97 1.38 1.64 ;
        RECT 1.23 0.97 1.38 1.44 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.88 1.2 7 1.44 ;
        RECT 6.45 1.315 7 1.435 ;
        RECT 6.45 1.175 6.6 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.48 0.885 8.63 1.145 ;
        RECT 8.38 1.025 8.5 1.385 ;
    END
  END SE
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.68 1.265 8.92 1.385 ;
        RECT 8.8 0.885 8.92 1.385 ;
        RECT 8.77 0.885 8.92 1.145 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.14 1.24 10.425 1.47 ;
        RECT 10.165 1.22 10.425 1.47 ;
    END
  END D1
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 0.94 10.715 1.09 ;
        RECT 10.545 0.94 10.665 1.18 ;
        RECT 9.86 0.97 10.715 1.09 ;
        RECT 9.4 1 10.045 1.12 ;
        RECT 9.28 1.265 9.52 1.385 ;
        RECT 9.4 1 9.52 1.385 ;
    END
  END S0
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 1.295 0.72 2.21 ;
        RECT 0.36 1.175 0.7 1.435 ;
        RECT 0.58 0.62 0.7 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.42 -0.18 10.54 0.82 ;
        RECT 9.14 -0.18 9.26 0.64 ;
        RECT 6.94 -0.18 7.06 0.79 ;
        RECT 4.75 0.49 4.99 0.61 ;
        RECT 4.87 -0.18 4.99 0.61 ;
        RECT 2.53 0.5 2.77 0.62 ;
        RECT 2.65 -0.18 2.77 0.62 ;
        RECT 0.94 0.49 1.18 0.61 ;
        RECT 0.94 -0.18 1.06 0.61 ;
        RECT 0.16 -0.18 0.28 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.22 1.83 10.34 2.79 ;
        RECT 8.84 1.745 8.96 2.79 ;
        RECT 6.8 1.85 6.92 2.79 ;
        RECT 4.71 2.01 4.95 2.13 ;
        RECT 4.71 2.01 4.83 2.79 ;
        RECT 2.49 1.88 2.73 2 ;
        RECT 2.49 1.88 2.61 2.79 ;
        RECT 1.02 1.56 1.14 2.79 ;
        RECT 0.18 1.56 0.3 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.96 0.82 10.955 0.82 10.955 1.71 10.82 1.71 10.82 1.83 10.7 1.83 10.7 1.71 9.72 1.71 9.72 1.24 9.84 1.24 9.84 1.59 10.835 1.59 10.835 0.7 10.84 0.7 10.84 0.58 10.96 0.58 ;
      POLYGON 9.9 0.85 9.74 0.85 9.74 0.88 9.16 0.88 9.16 1.505 9.6 1.505 9.6 2.21 9.48 2.21 9.48 1.625 8.26 1.625 8.26 1.68 8.04 1.68 8.04 2.01 7.92 2.01 7.92 1.56 8.14 1.56 8.14 0.77 8.12 0.77 8.12 0.65 8.36 0.65 8.36 0.77 8.26 0.77 8.26 1.505 9.04 1.505 9.04 0.76 9.62 0.76 9.62 0.73 9.78 0.73 9.78 0.59 9.9 0.59 ;
      POLYGON 8.74 0.765 8.62 0.765 8.62 0.53 8 0.53 8 0.89 8.02 0.89 8.02 1.44 7.8 1.44 7.8 2.13 8.36 2.13 8.36 1.865 8.48 1.865 8.48 2.25 7.68 2.25 7.68 1.44 7.36 1.44 7.36 1.2 7.48 1.2 7.48 1.32 7.9 1.32 7.9 1.01 7.88 1.01 7.88 0.41 8.74 0.41 ;
      POLYGON 7.76 0.77 7.64 0.77 7.64 1.03 7.24 1.03 7.24 1.56 7.56 1.56 7.56 2.21 7.44 2.21 7.44 1.68 6.19 1.68 6.19 1.82 6.07 1.82 6.07 1.47 6.13 1.47 6.13 0.72 6.07 0.72 6.07 0.6 6.31 0.6 6.31 0.72 6.25 0.72 6.25 1.56 7.12 1.56 7.12 0.91 7.52 0.91 7.52 0.65 7.76 0.65 ;
      POLYGON 6.64 0.79 6.52 0.79 6.52 0.48 5.95 0.48 5.95 1.11 6.01 1.11 6.01 1.35 5.95 1.35 5.95 1.94 6.44 1.94 6.44 2.03 6.56 2.03 6.56 2.15 6.32 2.15 6.32 2.06 5.83 2.06 5.83 0.48 5.35 0.48 5.35 0.88 5.47 0.88 5.47 1.12 5.23 1.12 5.23 0.85 4.51 0.85 4.51 0.48 4.03 0.48 4.03 0.94 4.15 0.94 4.15 1.06 3.91 1.06 3.91 0.36 4.63 0.36 4.63 0.73 5.23 0.73 5.23 0.36 6.64 0.36 ;
      POLYGON 5.71 1.99 5.59 1.99 5.59 1.36 4.63 1.36 4.63 1.33 4.51 1.33 4.51 1.21 4.75 1.21 4.75 1.24 5.59 1.24 5.59 0.72 5.47 0.72 5.47 0.6 5.71 0.6 ;
      POLYGON 5.51 2.25 5.07 2.25 5.07 1.89 4.395 1.89 4.395 2.23 3.12 2.23 3.12 1.76 1.62 1.76 1.62 1.8 1.5 1.8 1.5 1.56 1.54 1.56 1.54 0.68 1.78 0.68 1.78 0.8 1.66 0.8 1.66 1.64 3.12 1.64 3.12 1.1 3.03 1.1 3.03 0.98 3.27 0.98 3.27 1.1 3.24 1.1 3.24 2.11 3.65 2.11 3.65 1.13 3.77 1.13 3.77 2.11 4.275 2.11 4.275 1.77 5.19 1.77 5.19 2.13 5.51 2.13 ;
      POLYGON 5.11 1.09 4.39 1.09 4.39 1.65 4.15 1.65 4.15 1.53 4.27 1.53 4.27 0.72 4.15 0.72 4.15 0.6 4.39 0.6 4.39 0.97 5.11 0.97 ;
      POLYGON 3.53 1.99 3.41 1.99 3.41 0.78 3.08 0.78 3.08 0.86 2.55 0.86 2.55 1.21 2.43 1.21 2.43 0.74 2.96 0.74 2.96 0.66 3.41 0.66 3.41 0.54 3.53 0.54 ;
      POLYGON 2.87 1.45 2.29 1.45 2.29 1.52 2.01 1.52 2.01 1.4 2.17 1.4 2.17 0.56 1.42 0.56 1.42 0.85 1.06 0.85 1.06 1.12 0.82 1.12 0.82 0.73 1.3 0.73 1.3 0.44 2.29 0.44 2.29 1.33 2.75 1.33 2.75 1.13 2.87 1.13 ;
  END
END SMDFFHQX2

MACRO MX4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X1 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.945 1.005 1.185 1.22 ;
        RECT 0.885 0.94 1.145 1.18 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.345 1.26 3.585 1.45 ;
        RECT 3.205 1.165 3.465 1.38 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.705 1.27 4.825 1.54 ;
        RECT 4.505 1.42 4.825 1.54 ;
        RECT 4.365 1.52 4.625 1.67 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 1.52 5.205 1.67 ;
        RECT 5.065 1.25 5.185 1.67 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.245 1.005 6.505 1.16 ;
        RECT 6.105 0.94 6.365 1.125 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.685 1.23 6.945 1.38 ;
        RECT 5.925 1.31 6.825 1.43 ;
        RECT 6.045 1.31 6.165 2.17 ;
        RECT 4.605 2.05 6.165 2.17 ;
        RECT 4.245 2.13 4.725 2.25 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.365 1.34 0.485 1.99 ;
        RECT 0.29 0.59 0.41 1.46 ;
        RECT 0.07 0.885 0.41 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.305 0.46 6.545 0.58 ;
        RECT 6.425 -0.18 6.545 0.58 ;
        RECT 5.005 -0.18 5.125 0.86 ;
        RECT 3.605 0.53 3.845 0.65 ;
        RECT 3.605 -0.18 3.725 0.65 ;
        RECT 0.65 0.46 0.89 0.58 ;
        RECT 0.65 -0.18 0.77 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 6.485 1.71 6.605 2.79 ;
        RECT 4.845 2.29 5.085 2.79 ;
        RECT 3.365 2.02 3.485 2.79 ;
        RECT 0.785 1.34 0.905 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.185 1.67 7.025 1.67 7.025 1.83 6.905 1.83 6.905 1.55 7.065 1.55 7.065 0.86 6.845 0.86 6.845 0.82 6.065 0.82 6.065 0.56 5.445 0.56 5.445 1.31 5.565 1.31 5.565 1.43 5.325 1.43 5.325 1.13 4.585 1.13 4.585 1.3 4.065 1.3 4.065 1.42 3.945 1.42 3.945 1.18 4.445 1.18 4.445 1.01 5.325 1.01 5.325 0.44 5.745 0.44 5.745 0.36 5.985 0.36 5.985 0.44 6.185 0.44 6.185 0.7 6.845 0.7 6.845 0.62 6.965 0.62 6.965 0.74 7.185 0.74 ;
      POLYGON 5.845 0.8 5.805 0.8 5.805 1.93 4.485 1.93 4.485 2.01 3.605 2.01 3.605 1.9 2.81 1.9 2.81 1.22 2.93 1.22 2.93 0.86 2.81 0.86 2.81 0.6 2.93 0.6 2.93 0.74 3.05 0.74 3.05 1.34 2.93 1.34 2.93 1.78 3.725 1.78 3.725 1.89 4.365 1.89 4.365 1.81 5.685 1.81 5.685 0.8 5.605 0.8 5.605 0.68 5.845 0.68 ;
      POLYGON 4.485 0.89 3.825 0.89 3.825 1.54 4.125 1.54 4.125 1.65 4.245 1.65 4.245 1.77 4.005 1.77 4.005 1.66 3.705 1.66 3.705 0.89 3.365 0.89 3.365 0.48 2.09 0.48 2.09 1.64 1.85 1.64 1.85 1.52 1.97 1.52 1.97 0.36 3.485 0.36 3.485 0.77 4.365 0.77 4.365 0.62 4.485 0.62 ;
      POLYGON 2.81 1.1 2.69 1.1 2.69 2.12 1.265 2.12 1.265 1.46 1.305 1.46 1.305 0.77 1.25 0.77 1.25 0.65 1.49 0.65 1.49 0.77 1.425 0.77 1.425 1.58 1.385 1.58 1.385 2 2.57 2 2.57 0.98 2.81 0.98 ;
      POLYGON 2.51 0.84 2.45 0.84 2.45 1.88 1.61 1.88 1.61 0.53 1.13 0.53 1.13 0.82 0.765 0.82 0.765 1.15 0.645 1.15 0.645 0.7 1.01 0.7 1.01 0.41 1.73 0.41 1.73 1.76 2.33 1.76 2.33 0.72 2.39 0.72 2.39 0.6 2.51 0.6 ;
  END
END MX4X1

MACRO NOR3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 0.51 1.47 ;
        RECT 0.36 1 0.48 1.5 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.925 1.165 1.09 1.435 ;
        RECT 0.855 1.03 0.99 1.285 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.575 1 1.695 1.49 ;
        RECT 1.52 1 1.695 1.46 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.44 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.76 1.095 0.88 ;
        RECT 0.975 0.59 1.095 0.88 ;
        RECT 0.375 1.62 0.495 2.21 ;
        RECT 0.12 1.62 0.495 1.74 ;
        RECT 0.135 0.59 0.255 0.88 ;
        RECT 0.12 0.76 0.24 1.74 ;
        RECT 0.07 1.175 0.24 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.335 1.58 1.455 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 1.85 1.815 1.85 1.815 0.88 1.355 0.88 1.355 1.17 1.235 1.17 1.235 0.76 1.815 0.76 1.815 0.4 1.935 0.4 ;
  END
END NOR3BX1

MACRO INVXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVXL 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 1.04 0.24 1.455 ;
        RECT 0.07 1.04 0.24 1.445 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.68 0.675 1.695 ;
        RECT 0.36 1.175 0.675 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
        RECT 0.135 1.575 0.255 2.79 ;
    END
  END VDD
END INVXL

MACRO AND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X6 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 0.94 1.72 1.26 ;
        RECT 0.305 0.94 1.72 1.06 ;
        RECT 0.445 0.94 0.565 1.26 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.18 1.16 1.425 ;
        RECT 0.885 1.18 1.145 1.445 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 1.39 4.18 2.21 ;
        RECT 3.98 0.4 4.1 0.915 ;
        RECT 2.38 1.39 4.18 1.51 ;
        RECT 3.8 0.795 4.1 0.915 ;
        RECT 2.24 0.91 3.92 1.03 ;
        RECT 3.26 1.175 3.41 1.51 ;
        RECT 3.26 0.91 3.38 1.51 ;
        RECT 3.22 1.39 3.34 2.21 ;
        RECT 3.14 0.4 3.26 1.03 ;
        RECT 2.38 1.39 2.5 2.21 ;
        RECT 2.24 0.4 2.36 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.56 -0.18 3.68 0.79 ;
        RECT 2.72 -0.18 2.84 0.79 ;
        RECT 1.76 0.46 2 0.58 ;
        RECT 1.76 -0.18 1.88 0.58 ;
        RECT 0.48 -0.18 0.6 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.64 1.63 3.76 2.79 ;
        RECT 2.8 1.63 2.92 2.79 ;
        RECT 1.96 1.805 2.08 2.79 ;
        RECT 1.12 1.805 1.24 2.79 ;
        RECT 0.28 1.56 0.4 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.14 1.27 1.96 1.27 1.96 1.685 1.66 1.685 1.66 2.21 1.54 2.21 1.54 1.685 0.82 1.685 0.82 2.21 0.7 2.21 0.7 1.565 1.54 1.565 1.54 1.56 1.66 1.56 1.66 1.565 1.84 1.565 1.84 0.82 1.06 0.82 1.06 0.7 1.96 0.7 1.96 1.15 3.14 1.15 ;
  END
END AND2X6

MACRO SEDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX8 0 0 ;
  SIZE 14.79 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 1.465 2.775 2.21 ;
        RECT 2.655 0.68 2.775 1.005 ;
        RECT 2.635 0.885 2.755 1.585 ;
        RECT 0.07 1.005 2.755 1.125 ;
        RECT 1.815 0.68 1.935 2.21 ;
        RECT 0.975 0.68 1.095 2.205 ;
        RECT 0.135 0.68 0.255 2.205 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 1.15 5.15 1.47 ;
        RECT 4.91 1.15 5.15 1.465 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.305 1.22 10.665 1.35 ;
        RECT 10.165 1.23 10.425 1.395 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.25 1.14 12.4 1.61 ;
        RECT 12.255 1.14 12.375 1.64 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.935 1.21 14.195 1.465 ;
        RECT 13.855 1.21 14.195 1.44 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.315 0.97 14.435 1.21 ;
        RECT 13.135 0.97 14.435 1.09 ;
        RECT 13.615 0.94 13.905 1.09 ;
        RECT 13.615 0.92 13.735 1.16 ;
        RECT 13.135 0.97 13.255 1.26 ;
        RECT 13.055 1.14 13.175 1.44 ;
    END
  END E
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.79 0.18 ;
        RECT 14.115 -0.18 14.235 0.82 ;
        RECT 12.535 0.6 12.775 0.72 ;
        RECT 12.535 -0.18 12.655 0.72 ;
        RECT 10.465 -0.18 10.585 0.65 ;
        RECT 9.505 -0.18 9.625 0.63 ;
        RECT 7.07 0.5 7.31 0.62 ;
        RECT 7.07 -0.18 7.19 0.62 ;
        RECT 5.37 0.43 5.61 0.55 ;
        RECT 5.49 -0.18 5.61 0.55 ;
        RECT 3.915 -0.18 4.035 0.67 ;
        RECT 3.075 -0.18 3.195 0.67 ;
        RECT 2.235 -0.18 2.355 0.67 ;
        RECT 1.395 -0.18 1.515 0.67 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.79 2.79 ;
        RECT 13.935 1.825 14.055 2.79 ;
        RECT 12.455 2.28 12.695 2.79 ;
        RECT 10.345 1.94 10.585 2.09 ;
        RECT 10.345 1.94 10.465 2.79 ;
        RECT 9.505 2.14 9.625 2.79 ;
        RECT 7.43 1.94 7.67 2.06 ;
        RECT 7.43 1.94 7.55 2.79 ;
        RECT 5.07 2.11 5.19 2.79 ;
        RECT 3.915 1.56 4.035 2.79 ;
        RECT 3.075 1.56 3.195 2.79 ;
        RECT 2.235 1.465 2.355 2.79 ;
        RECT 1.395 1.465 1.515 2.79 ;
        RECT 0.555 1.465 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.675 1.705 14.535 1.705 14.535 1.825 14.415 1.825 14.415 1.705 13.615 1.705 13.615 1.42 13.375 1.42 13.375 1.3 13.735 1.3 13.735 1.585 14.555 1.585 14.555 0.85 14.535 0.85 14.535 0.58 14.655 0.58 14.655 0.73 14.675 0.73 ;
      POLYGON 13.595 0.8 13.015 0.8 13.015 1.02 12.935 1.02 12.935 1.56 13.335 1.56 13.335 2.21 13.215 2.21 13.215 1.68 12.815 1.68 12.815 1.02 12.005 1.02 12.005 1.44 11.855 1.44 11.855 1.68 11.585 1.68 11.585 1.56 11.735 1.56 11.735 1.32 11.885 1.32 11.885 0.84 11.785 0.84 11.785 0.6 11.905 0.6 11.905 0.72 12.005 0.72 12.005 0.9 12.895 0.9 12.895 0.68 13.475 0.68 13.475 0.56 13.595 0.56 ;
      POLYGON 12.695 2.12 12.43 2.12 12.43 2.16 12.165 2.16 12.165 2.25 10.72 2.25 10.72 1.82 10.105 1.82 10.105 2.15 9.985 2.15 9.985 1.635 9.925 1.635 9.925 0.99 9.985 0.99 9.985 0.6 10.105 0.6 10.105 1.11 10.045 1.11 10.045 1.515 10.105 1.515 10.105 1.7 10.84 1.7 10.84 2.13 12.045 2.13 12.045 2.04 12.31 2.04 12.31 2 12.575 2 12.575 1.22 12.695 1.22 ;
      POLYGON 12.295 0.78 12.175 0.78 12.175 0.48 11.615 0.48 11.615 0.96 11.765 0.96 11.765 1.2 11.615 1.2 11.615 1.34 11.465 1.34 11.465 1.8 11.975 1.8 11.975 1.76 12.215 1.76 12.215 1.88 12.095 1.88 12.095 1.92 11.345 1.92 11.345 1.34 11.025 1.34 11.025 1.22 11.495 1.22 11.495 0.36 12.295 0.36 ;
      POLYGON 11.375 0.89 10.905 0.89 10.905 1.46 11.105 1.46 11.105 1.56 11.225 1.56 11.225 2.01 10.985 2.01 10.985 1.58 10.785 1.58 10.785 0.89 10.225 0.89 10.225 0.48 9.865 0.48 9.865 0.87 9.265 0.87 9.265 0.54 8.31 0.54 8.31 0.91 8.87 0.91 8.87 1.77 8.75 1.77 8.75 1.03 8.19 1.03 8.19 0.42 9.385 0.42 9.385 0.75 9.745 0.75 9.745 0.36 10.345 0.36 10.345 0.77 11.255 0.77 11.255 0.6 11.375 0.6 ;
      POLYGON 9.805 1.52 9.65 1.52 9.65 2.02 9.385 2.02 9.385 2.25 7.79 2.25 7.79 1.82 7.31 1.82 7.31 2.25 5.335 2.25 5.335 1.99 4.455 1.99 4.455 2.21 4.335 2.21 4.335 1.44 3.615 1.44 3.615 2.21 3.495 2.21 3.495 1.245 2.875 1.245 2.875 1.125 3.495 1.125 3.495 0.62 3.615 0.62 3.615 1.32 4.395 1.32 4.395 0.62 4.515 0.62 4.515 1.44 4.455 1.44 4.455 1.87 5.27 1.87 5.27 1.15 5.39 1.15 5.39 1.87 5.455 1.87 5.455 2.13 7.19 2.13 7.19 1.7 7.91 1.7 7.91 2.13 9.265 2.13 9.265 1.9 9.53 1.9 9.53 1.4 9.685 1.4 9.685 1.16 9.805 1.16 ;
      POLYGON 9.26 1.78 9.145 1.78 9.145 2.01 8.03 2.01 8.03 1.58 7.07 1.58 7.07 2.01 5.63 2.01 5.63 1.15 5.75 1.15 5.75 1.89 6.47 1.89 6.47 0.86 6.59 0.86 6.59 1.89 6.95 1.89 6.95 1.46 7.71 1.46 7.71 1.1 7.59 1.1 7.59 0.98 7.83 0.98 7.83 1.46 8.15 1.46 8.15 1.89 8.51 1.89 8.51 1.15 8.63 1.15 8.63 1.89 9.025 1.89 9.025 0.78 8.905 0.78 8.905 0.66 9.145 0.66 9.145 1.5 9.26 1.5 ;
      POLYGON 8.39 1.77 8.27 1.77 8.27 1.34 7.95 1.34 7.95 0.78 7.55 0.78 7.55 0.86 7.07 0.86 7.07 1.1 6.95 1.1 6.95 0.74 7.43 0.74 7.43 0.66 7.77 0.66 7.77 0.54 7.89 0.54 7.89 0.66 8.07 0.66 8.07 1.22 8.39 1.22 ;
      POLYGON 7.47 1.31 7.35 1.31 7.35 1.34 6.83 1.34 6.83 1.77 6.71 1.77 6.71 0.54 6.83 0.54 6.83 1.22 7.23 1.22 7.23 1.19 7.47 1.19 ;
      POLYGON 6.35 1.77 6.23 1.77 6.23 0.78 6.045 0.78 6.045 0.79 5.13 0.79 5.13 0.48 4.275 0.48 4.275 1.2 4.155 1.2 4.155 0.36 5.25 0.36 5.25 0.67 5.925 0.67 5.925 0.66 6.23 0.66 6.23 0.54 6.35 0.54 ;
      POLYGON 6.11 1.15 5.99 1.15 5.99 1.03 4.79 1.03 4.79 1.59 4.765 1.59 4.765 1.71 4.645 1.71 4.645 1.47 4.67 1.47 4.67 0.6 5.01 0.6 5.01 0.72 4.79 0.72 4.79 0.91 6.11 0.91 ;
  END
END SEDFFHQX8

MACRO DFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX2 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.885 0.415 1.37 ;
        RECT 0.07 0.885 0.415 1.34 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.07 1.09 1.435 ;
        RECT 0.835 0.915 0.955 1.29 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.79 1.005 6.03 1.18 ;
        RECT 5.87 0.8 6.02 1.18 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.61 1.36 6.73 2.01 ;
        RECT 6.57 0.74 6.69 1.48 ;
        RECT 6.45 0.74 6.69 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.41 0.74 7.65 0.86 ;
        RECT 7.45 1.3 7.57 2.01 ;
        RECT 7.41 0.74 7.53 1.42 ;
        RECT 7.32 0.885 7.53 1.145 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.95 -0.18 8.07 0.38 ;
        RECT 6.93 -0.18 7.17 0.38 ;
        RECT 5.97 -0.18 6.21 0.38 ;
        RECT 4.74 -0.18 4.86 0.76 ;
        RECT 2.96 0.35 3.2 0.47 ;
        RECT 2.96 -0.18 3.08 0.47 ;
        RECT 0.91 -0.18 1.03 0.75 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.87 1.36 7.99 2.79 ;
        RECT 7.03 1.36 7.15 2.79 ;
        RECT 6.19 1.36 6.31 2.79 ;
        RECT 4.78 2.16 5.02 2.28 ;
        RECT 4.78 2.16 4.9 2.79 ;
        RECT 2.98 2.23 3.22 2.79 ;
        RECT 1.035 2.01 1.155 2.79 ;
        RECT 0.135 1.49 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.55 1.18 8.47 1.18 8.47 1.6 8.35 1.6 8.35 1.18 7.67 1.18 7.67 1.06 8.43 1.06 8.43 0.68 8.55 0.68 ;
      POLYGON 8.45 0.52 8.31 0.52 8.31 0.62 6.985 0.62 6.985 1.24 6.865 1.24 6.865 0.62 6.33 0.62 6.33 1.24 6.21 1.24 6.21 0.62 5.28 0.62 5.28 0.76 5.3 0.76 5.3 1.68 5.5 1.68 5.5 1.8 5.18 1.8 5.18 1.52 4.82 1.52 4.82 1.28 4.94 1.28 4.94 1.4 5.18 1.4 5.18 0.88 5.16 0.88 5.16 0.5 8.19 0.5 8.19 0.4 8.45 0.4 ;
      POLYGON 5.83 2.04 4.515 2.04 4.515 2.11 4.105 2.11 4.105 2.25 3.865 2.25 3.865 2.11 2.66 2.11 2.66 2.25 2.42 2.25 2.42 2.13 2.54 2.13 2.54 1.99 4.395 1.99 4.395 1.92 5.71 1.92 5.71 1.48 5.55 1.48 5.55 0.86 5.49 0.86 5.49 0.74 5.73 0.74 5.73 0.86 5.67 0.86 5.67 1.36 5.83 1.36 ;
      POLYGON 5.06 1.12 4.7 1.12 4.7 1.73 4.26 1.73 4.26 1.87 4.14 1.87 4.14 1.61 4.58 1.61 4.58 1.12 4.04 1.12 4.04 0.62 4.16 0.62 4.16 1 5.06 1 ;
      POLYGON 4.46 1.49 3.8 1.49 3.8 1.31 3.72 1.31 3.72 1.07 3.8 1.07 3.8 0.5 3.44 0.5 3.44 0.71 2.72 0.71 2.72 0.5 2.11 0.5 2.11 1.37 2.2 1.37 2.2 1.49 1.96 1.49 1.96 1.37 1.99 1.37 1.99 0.5 1.58 0.5 1.58 0.51 1.45 0.51 1.45 1.37 1.6 1.37 1.6 1.61 1.48 1.61 1.48 1.49 1.33 1.49 1.33 0.39 1.46 0.39 1.46 0.38 2.4 0.38 2.4 0.36 2.64 0.36 2.64 0.38 2.84 0.38 2.84 0.59 3.32 0.59 3.32 0.38 3.92 0.38 3.92 1.37 4.46 1.37 ;
      POLYGON 3.68 0.95 3.6 0.95 3.6 1.63 3.64 1.63 3.64 1.87 3.52 1.87 3.52 1.75 3.48 1.75 3.48 1.49 2.78 1.49 2.78 1.37 3.48 1.37 3.48 0.83 3.56 0.83 3.56 0.62 3.68 0.62 ;
      POLYGON 3.36 1.25 2.46 1.25 2.46 1.87 2.34 1.87 2.34 0.8 2.26 0.8 2.26 0.68 2.5 0.68 2.5 0.8 2.46 0.8 2.46 1.13 3.36 1.13 ;
      POLYGON 2.04 1.87 1.92 1.87 1.92 1.85 0.555 1.85 0.555 1.61 0.535 1.61 0.535 0.765 0.27 0.765 0.27 0.51 0.39 0.51 0.39 0.645 0.655 0.645 0.655 1.49 0.675 1.49 0.675 1.73 1.72 1.73 1.72 0.62 1.84 0.62 1.84 1.63 2.04 1.63 ;
  END
END DFFTRX2

MACRO TLATNTSCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX4 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.705 0.59 6.825 2.21 ;
        RECT 5.87 1.025 6.825 1.145 ;
        RECT 5.865 0.885 6.02 1.025 ;
        RECT 5.885 0.885 6.005 1.68 ;
        RECT 5.865 1.56 5.985 2.21 ;
        RECT 5.865 0.59 5.985 1.025 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.175 0.435 1.295 ;
        RECT 0.315 1.055 0.435 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.165 1.145 1.4 ;
        RECT 0.795 1.165 1.145 1.375 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 1.52 1.435 1.755 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 7.125 -0.18 7.245 0.64 ;
        RECT 6.285 -0.18 6.405 0.64 ;
        RECT 5.445 -0.18 5.565 0.64 ;
        RECT 4.415 -0.18 4.535 0.9 ;
        RECT 3.065 0.68 3.305 0.8 ;
        RECT 3.185 -0.18 3.305 0.8 ;
        RECT 0.955 0.685 1.195 0.805 ;
        RECT 0.955 -0.18 1.075 0.805 ;
        RECT 0.175 -0.18 0.295 0.865 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 7.125 1.56 7.245 2.79 ;
        RECT 6.285 1.56 6.405 2.79 ;
        RECT 5.445 1.6 5.565 2.79 ;
        RECT 4.625 1.8 4.745 2.79 ;
        RECT 4.605 1.56 4.725 1.92 ;
        RECT 3.255 2.29 3.495 2.79 ;
        RECT 1.015 1.9 1.135 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.765 1.385 5.445 1.385 5.445 1.48 5.145 1.48 5.145 2.21 5.025 2.21 5.025 1.36 5.325 1.36 5.325 0.88 5.055 0.88 5.055 0.64 5.175 0.64 5.175 0.76 5.445 0.76 5.445 1.265 5.765 1.265 ;
      POLYGON 5.205 1.24 5.085 1.24 5.085 1.14 4.175 1.14 4.175 0.54 3.765 0.54 3.765 0.74 3.815 0.74 3.815 1.57 3.975 1.57 3.975 1.69 3.695 1.69 3.695 1.04 2.825 1.04 2.825 0.56 2.305 0.56 2.305 1.64 2.185 1.64 2.185 0.44 2.565 0.44 2.565 0.36 2.805 0.36 2.805 0.44 2.945 0.44 2.945 0.92 3.545 0.92 3.545 0.62 3.645 0.62 3.645 0.42 4.295 0.42 4.295 1.02 5.085 1.02 5.085 1 5.205 1 ;
      POLYGON 4.865 1.42 4.305 1.42 4.305 1.93 3.145 1.93 3.145 1.6 3.025 1.6 3.025 1.48 3.265 1.48 3.265 1.81 4.185 1.81 4.185 1.38 3.935 1.38 3.935 0.66 4.055 0.66 4.055 1.26 4.305 1.26 4.305 1.3 4.865 1.3 ;
      POLYGON 4.505 2.18 4 2.18 4 2.17 2.425 2.17 2.425 0.68 2.665 0.68 2.665 0.8 2.545 0.8 2.545 1.86 2.705 1.86 2.705 2.05 4.12 2.05 4.12 2.06 4.505 2.06 ;
      POLYGON 3.485 1.28 3.365 1.28 3.365 1.34 2.665 1.34 2.665 1.22 3.245 1.22 3.245 1.16 3.485 1.16 ;
      POLYGON 2.285 2 2.165 2 2.165 1.88 1.945 1.88 1.945 0.505 1.435 0.505 1.435 1.045 0.675 1.045 0.675 1.96 0.315 1.96 0.315 1.84 0.555 1.84 0.555 0.805 0.595 0.805 0.595 0.625 0.715 0.625 0.715 0.925 1.315 0.925 1.315 0.385 2.065 0.385 2.065 1.76 2.285 1.76 ;
      POLYGON 1.825 1.4 1.675 1.4 1.675 1.995 1.555 1.995 1.555 2.115 1.435 2.115 1.435 1.875 1.555 1.875 1.555 0.625 1.675 0.625 1.675 1.16 1.825 1.16 ;
  END
END TLATNTSCAX4

MACRO DFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX4 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.995 0.72 2.235 0.84 ;
        RECT 2.075 1.28 2.195 2.11 ;
        RECT 2.035 0.72 2.155 1.4 ;
        RECT 1.23 1.025 2.155 1.145 ;
        RECT 1.23 0.885 1.38 1.145 ;
        RECT 1.235 0.72 1.355 2.11 ;
        RECT 1.23 0.72 1.355 1.145 ;
        RECT 1.035 0.72 1.355 0.84 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.06 0.51 1.435 ;
        RECT 0.375 0.84 0.495 1.435 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.395 1.23 6.655 1.46 ;
        RECT 6.455 1.1 6.575 1.51 ;
    END
  END D
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.675 -0.18 6.795 0.74 ;
        RECT 5.095 -0.18 5.335 0.36 ;
        RECT 3.555 -0.18 3.675 0.38 ;
        RECT 2.475 -0.18 2.715 0.36 ;
        RECT 1.515 -0.18 1.755 0.36 ;
        RECT 0.555 -0.18 0.675 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.575 1.87 6.695 2.79 ;
        RECT 4.995 2.29 5.235 2.79 ;
        RECT 3.335 1.75 3.455 2.79 ;
        RECT 2.495 1.59 2.615 2.79 ;
        RECT 1.655 1.46 1.775 2.79 ;
        RECT 0.815 1.46 0.935 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.335 0.84 7.255 0.84 7.255 1.42 7.115 1.42 7.115 1.99 6.995 1.99 6.995 1.75 6.195 1.75 6.195 2.17 4.275 2.17 4.275 1.65 3.975 1.65 3.975 1.41 4.095 1.41 4.095 1.53 4.515 1.53 4.515 1 4.635 1 4.635 1.65 4.395 1.65 4.395 2.05 6.075 2.05 6.075 1.43 6.195 1.43 6.195 1.63 6.995 1.63 6.995 1.3 7.135 1.3 7.135 0.84 7.095 0.84 7.095 0.72 7.335 0.72 ;
      POLYGON 7.015 1.18 6.775 1.18 6.775 0.98 6.255 0.98 6.255 1.24 6.135 1.24 6.135 0.54 5.725 0.54 5.725 0.6 5.715 0.6 5.715 1.65 5.595 1.65 5.595 0.6 4.81 0.6 4.81 0.54 4.115 0.54 4.115 0.62 3.315 0.62 3.315 0.6 0.915 0.6 0.915 0.66 0.255 0.66 0.255 0.9 0.24 0.9 0.24 1.555 0.515 1.555 0.515 1.795 0.395 1.795 0.395 1.675 0.12 1.675 0.12 0.78 0.135 0.78 0.135 0.54 0.795 0.54 0.795 0.48 3.435 0.48 3.435 0.5 3.995 0.5 3.995 0.4 4.235 0.4 4.235 0.42 4.93 0.42 4.93 0.48 5.605 0.48 5.605 0.42 6.255 0.42 6.255 0.86 6.895 0.86 6.895 1.06 7.015 1.06 ;
      POLYGON 6.015 1.31 5.955 1.31 5.955 1.93 5.715 1.93 5.715 1.89 5.355 1.89 5.355 1.59 4.995 1.59 4.995 1.47 5.475 1.47 5.475 1.77 5.835 1.77 5.835 1.19 5.895 1.19 5.895 0.66 6.015 0.66 ;
      POLYGON 5.395 1.29 4.875 1.29 4.875 1.93 4.515 1.93 4.515 1.81 4.755 1.81 4.755 0.84 4.615 0.84 4.615 0.72 4.875 0.72 4.875 1.17 5.275 1.17 5.275 1.05 5.395 1.05 ;
      POLYGON 4.375 1.29 3.855 1.29 3.855 1.77 4.035 1.77 4.035 1.81 4.155 1.81 4.155 1.93 3.915 1.93 3.915 1.89 3.735 1.89 3.735 1.49 3.175 1.49 3.175 1.25 3.295 1.25 3.295 1.37 3.735 1.37 3.735 1.17 4.255 1.17 4.255 0.66 4.375 0.66 ;
      POLYGON 3.615 1.25 3.495 1.25 3.495 1.13 3.035 1.13 3.035 2.11 2.915 2.11 2.915 1.13 2.515 1.13 2.515 1.16 2.275 1.16 2.275 1.01 3.075 1.01 3.075 0.84 2.955 0.84 2.955 0.72 3.195 0.72 3.195 1.01 3.615 1.01 ;
  END
END DFFQX4

MACRO AND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X8 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.42 0.75 2.54 1.22 ;
        RECT 0.39 0.75 2.54 0.87 ;
        RECT 0.42 0.75 0.54 1.22 ;
        RECT 0.36 0.885 0.54 1.145 ;
        RECT 0.39 0.75 0.54 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.175 2.25 1.435 ;
        RECT 2.1 0.99 2.22 1.435 ;
        RECT 1.225 0.99 2.22 1.11 ;
        RECT 0.98 1.04 1.345 1.16 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.23 1.725 1.5 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.64 0.715 5.88 0.835 ;
        RECT 5.72 1.295 5.84 2.21 ;
        RECT 3.18 0.765 5.76 0.885 ;
        RECT 3.2 1.295 5.84 1.415 ;
        RECT 4.9 0.765 5.15 1.145 ;
        RECT 4.8 0.715 5.04 0.885 ;
        RECT 4.9 0.715 5.02 1.415 ;
        RECT 4.88 1.295 5 2.21 ;
        RECT 3.96 0.715 4.2 0.885 ;
        RECT 4.04 1.295 4.16 2.21 ;
        RECT 3.2 1.295 3.32 2.21 ;
        RECT 3.06 0.715 3.3 0.835 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.28 -0.18 5.4 0.645 ;
        RECT 4.44 -0.18 4.56 0.645 ;
        RECT 3.54 -0.18 3.66 0.64 ;
        RECT 2.58 -0.18 2.82 0.39 ;
        RECT 0.5 0.51 0.74 0.63 ;
        RECT 0.5 -0.18 0.62 0.63 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.3 1.535 5.42 2.79 ;
        RECT 4.46 1.535 4.58 2.79 ;
        RECT 3.62 1.535 3.74 2.79 ;
        RECT 2.78 1.86 2.9 2.79 ;
        RECT 1.94 1.86 2.06 2.79 ;
        RECT 1.1 1.86 1.22 2.79 ;
        RECT 0.26 1.56 0.38 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.78 1.175 2.78 1.175 2.78 1.74 2.48 1.74 2.48 2.21 2.36 2.21 2.36 1.74 1.64 1.74 1.64 2.21 1.52 2.21 1.52 1.74 0.8 1.74 0.8 2.21 0.68 2.21 0.68 1.56 0.8 1.56 0.8 1.62 2.36 1.62 2.36 1.56 2.48 1.56 2.48 1.62 2.66 1.62 2.66 0.63 1.56 0.63 1.56 0.51 2.78 0.51 2.78 1.055 4.78 1.055 ;
  END
END AND3X8

MACRO AOI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X1 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.04 1.09 1.16 ;
        RECT 0.94 0.885 1.09 1.16 ;
        RECT 0.815 1.04 0.935 1.295 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.295 2.48 1.425 ;
        RECT 2.1 1.15 2.25 1.435 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.77 0.51 1.145 ;
        RECT 0.36 0.77 0.48 1.38 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.94 1.98 1.4 ;
        RECT 1.81 1 1.96 1.435 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.965 1.67 1.435 ;
        RECT 1.54 0.94 1.66 1.44 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6141 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.64 0.82 2.76 2.205 ;
        RECT 2.42 0.82 2.76 0.94 ;
        RECT 1.44 0.7 2.56 0.82 ;
        RECT 2.44 0.58 2.56 0.94 ;
        RECT 2.39 0.595 2.56 0.855 ;
        RECT 1.32 0.65 1.56 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.96 0.46 2.2 0.58 ;
        RECT 1.96 -0.18 2.08 0.58 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.035 2.19 1.155 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.34 2.25 1.38 2.25 1.38 1.8 1.5 1.8 1.5 2.13 2.22 2.13 2.22 1.555 2.34 1.555 ;
      POLYGON 1.92 2.01 1.8 2.01 1.8 1.68 0.675 1.68 0.675 2.21 0.555 2.21 0.555 1.56 1.8 1.56 1.8 1.555 1.92 1.555 ;
  END
END AOI221X1

MACRO TLATNX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX2 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.465 0.94 5.785 1.09 ;
        RECT 5.465 0.64 5.585 1.99 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 0.885 3.99 1.145 ;
        RECT 3.785 0.64 3.905 1.99 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 0.94 3.175 1.21 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.07 0.875 1.19 ;
        RECT 0.305 1.23 0.715 1.38 ;
        RECT 0.595 1.07 0.715 1.38 ;
    END
  END D
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.885 1.34 6.005 2.79 ;
        RECT 5.045 1.34 5.165 2.79 ;
        RECT 4.205 1.34 4.325 2.79 ;
        RECT 3.305 1.4 3.545 1.64 ;
        RECT 3.305 1.4 3.425 2.79 ;
        RECT 2.055 2.27 2.295 2.79 ;
        RECT 0.735 1.81 0.855 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.885 -0.18 6.005 0.69 ;
        RECT 5.045 -0.18 5.165 0.69 ;
        RECT 4.205 -0.18 4.325 0.69 ;
        RECT 3.245 -0.18 3.485 0.34 ;
        RECT 2.015 -0.18 2.135 0.71 ;
        RECT 0.555 -0.18 0.675 0.71 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.345 1.2 4.745 1.2 4.745 1.99 4.625 1.99 4.625 0.64 4.745 0.64 4.745 1.08 5.345 1.08 ;
      POLYGON 3.625 1.2 3.505 1.2 3.505 0.82 3.23 0.82 3.23 0.58 2.555 0.58 2.555 1.79 2.775 1.79 2.775 1.91 2.435 1.91 2.435 1.43 2.175 1.43 2.175 1.55 2.055 1.55 2.055 1.31 2.435 1.31 2.435 0.46 3.35 0.46 3.35 0.7 3.625 0.7 ;
      POLYGON 3.065 2.15 1.115 2.15 1.115 1.55 1.535 1.55 1.535 1.07 1.035 1.07 1.035 0.95 0.475 0.95 0.475 1.07 0.355 1.07 0.355 0.83 1.655 0.83 1.655 1.35 1.695 1.35 1.695 1.59 1.655 1.59 1.655 1.67 1.235 1.67 1.235 2.03 2.945 2.03 2.945 1.46 2.675 1.46 2.675 0.7 3.005 0.7 3.005 0.82 2.795 0.82 2.795 1.34 3.065 1.34 ;
      POLYGON 2.315 1.15 1.935 1.15 1.935 1.91 1.355 1.91 1.355 1.79 1.815 1.79 1.815 1.15 1.775 1.15 1.775 0.71 1.195 0.71 1.195 0.47 1.315 0.47 1.315 0.59 1.895 0.59 1.895 1.03 2.315 1.03 ;
      POLYGON 1.415 1.43 0.955 1.43 0.955 1.62 0.435 1.62 0.435 1.93 0.315 1.93 0.315 1.74 0.065 1.74 0.065 0.59 0.135 0.59 0.135 0.47 0.255 0.47 0.255 0.71 0.185 0.71 0.185 1.5 0.835 1.5 0.835 1.31 1.415 1.31 ;
  END
END TLATNX2

MACRO SDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX1 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 1.22 2.25 1.46 ;
        RECT 1.755 1.52 2.15 1.67 ;
        RECT 2.03 1.34 2.15 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.915 1.29 7.035 1.53 ;
        RECT 6.74 1.29 7.035 1.435 ;
        RECT 6.74 1.175 6.89 1.435 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.115 1.23 8.395 1.47 ;
        RECT 8.135 1.21 8.395 1.47 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 0.94 8.685 1.09 ;
        RECT 8.475 0.85 8.595 1.09 ;
        RECT 7.515 0.95 8.685 1.07 ;
        RECT 7.755 0.87 7.995 1.07 ;
        RECT 7.395 1.41 7.635 1.53 ;
        RECT 7.515 0.95 7.635 1.53 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.885 1.67 1.145 ;
        RECT 1.455 0.885 1.575 2.21 ;
        RECT 1.395 0.68 1.515 1.025 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.315 -0.18 8.435 0.73 ;
        RECT 7.035 -0.18 7.155 0.73 ;
        RECT 4.845 -0.18 5.085 0.32 ;
        RECT 3.225 -0.18 3.465 0.32 ;
        RECT 1.755 0.55 1.995 0.67 ;
        RECT 1.755 -0.18 1.875 0.67 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 8.315 1.83 8.435 2.79 ;
        RECT 6.835 1.89 7.075 2.01 ;
        RECT 6.835 1.89 6.955 2.79 ;
        RECT 4.865 2.16 4.985 2.79 ;
        RECT 3.205 2.16 3.445 2.28 ;
        RECT 3.205 2.16 3.325 2.79 ;
        RECT 1.875 1.79 1.995 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.925 1.83 8.855 1.83 8.855 1.95 8.735 1.95 8.735 1.71 7.875 1.71 7.875 1.31 7.755 1.31 7.755 1.19 7.995 1.19 7.995 1.59 8.805 1.59 8.805 0.82 8.735 0.82 8.735 0.49 8.855 0.49 8.855 0.7 8.925 0.7 ;
      POLYGON 7.795 0.75 7.395 0.75 7.395 1.29 7.275 1.29 7.275 1.65 7.655 1.65 7.655 1.95 7.535 1.95 7.535 1.77 6.165 1.77 6.165 1.88 6.045 1.88 6.045 1.64 6.145 1.64 6.145 0.66 6.265 0.66 6.265 1.65 7.155 1.65 7.155 1.17 7.275 1.17 7.275 0.63 7.675 0.63 7.675 0.49 7.795 0.49 ;
      POLYGON 6.795 0.67 6.555 0.67 6.555 0.54 6.025 0.54 6.025 1.08 5.925 1.08 5.925 1.28 6.005 1.28 6.005 1.52 5.925 1.52 5.925 2 6.375 2 6.375 1.89 6.615 1.89 6.615 2.01 6.495 2.01 6.495 2.12 5.805 2.12 5.805 0.96 5.905 0.96 5.905 0.54 5.38 0.54 5.38 0.56 4.325 0.56 4.325 1.22 4.205 1.22 4.205 0.44 5.26 0.44 5.26 0.42 5.405 0.42 5.405 0.4 5.645 0.4 5.645 0.42 6.675 0.42 6.675 0.55 6.795 0.55 ;
      POLYGON 5.785 0.84 5.685 0.84 5.685 1.86 5.565 1.86 5.565 1.48 4.725 1.48 4.725 1.36 5.565 1.36 5.565 0.84 5.545 0.84 5.545 0.72 5.785 0.72 ;
      POLYGON 5.605 2.24 5.325 2.24 5.325 2.04 4.595 2.04 4.595 2.1 4.425 2.1 4.425 2.24 4.185 2.24 4.185 2.1 3.68 2.1 3.68 2.04 2.355 2.04 2.355 1.68 2.37 1.68 2.37 1.1 2.355 1.1 2.355 0.68 2.475 0.68 2.475 0.98 2.49 0.98 2.49 1.8 2.475 1.8 2.475 1.92 3.68 1.92 3.68 1.16 3.605 1.16 3.605 1.04 3.845 1.04 3.845 1.16 3.8 1.16 3.8 1.98 4.475 1.98 4.475 1.92 5.445 1.92 5.445 2.12 5.605 2.12 ;
      POLYGON 5.185 1.22 4.565 1.22 4.565 1.8 4.325 1.8 4.325 1.68 4.445 1.68 4.445 0.72 4.685 0.72 4.685 0.84 4.565 0.84 4.565 1.1 5.065 1.1 5.065 0.98 5.185 0.98 ;
      POLYGON 4.085 1.86 3.965 1.86 3.965 0.9 3.925 0.9 3.925 0.66 2.985 0.66 2.985 0.5 2.845 0.5 2.845 0.38 3.105 0.38 3.105 0.54 4.045 0.54 4.045 0.78 4.085 0.78 ;
      POLYGON 3.485 1.24 2.865 1.24 2.865 1.68 2.965 1.68 2.965 1.8 2.725 1.8 2.725 1.68 2.745 1.68 2.745 0.78 2.605 0.78 2.605 0.56 2.235 0.56 2.235 0.91 1.91 0.91 1.91 1.24 1.79 1.24 1.79 0.79 2.115 0.79 2.115 0.44 2.725 0.44 2.725 0.66 2.865 0.66 2.865 1.12 3.485 1.12 ;
      POLYGON 1.155 1.58 1.035 1.58 1.035 1.32 1.005 1.32 1.005 1.2 0.375 1.2 0.375 1.08 1.005 1.08 1.005 0.68 1.125 0.68 1.125 1.2 1.155 1.2 ;
  END
END SDFFX1

MACRO ADDFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFXL 0 0 ;
  SIZE 7.54 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.78 5.97 0.9 ;
        RECT 2.625 0.72 3.355 0.8 ;
        RECT 2.705 0.78 5.97 0.84 ;
        RECT 2.625 0.65 2.885 0.8 ;
        RECT 2.705 0.65 2.825 0.96 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.49 1.02 6.61 1.5 ;
        RECT 6.45 1.02 6.61 1.435 ;
        RECT 2.045 1.08 6.61 1.14 ;
        RECT 3.585 1.02 6.61 1.14 ;
        RECT 2.26 1.08 3.705 1.2 ;
        RECT 1.445 1.02 2.38 1.08 ;
        RECT 1.445 0.96 2.165 1.08 ;
        RECT 1.325 1.08 1.565 1.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.975 1.26 6.33 1.38 ;
        RECT 1.805 1.32 4.095 1.44 ;
        RECT 2.915 1.32 3.175 1.67 ;
        RECT 1.805 1.2 1.925 1.44 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.605 0.675 1.965 ;
        RECT 0.155 1.005 0.675 1.125 ;
        RECT 0.555 0.645 0.675 1.125 ;
        RECT 0.07 1.605 0.675 1.725 ;
        RECT 0.07 1.465 0.275 1.725 ;
        RECT 0.155 1.005 0.275 1.725 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.175 0.4 7.295 0.64 ;
        RECT 7.03 1.465 7.18 1.725 ;
        RECT 7.055 0.52 7.175 1.725 ;
        RECT 7.05 1.465 7.17 2.09 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.54 0.18 ;
        RECT 6.755 -0.18 6.875 0.64 ;
        RECT 4.545 0.3 4.785 0.42 ;
        RECT 4.545 -0.18 4.665 0.42 ;
        RECT 3.705 -0.18 3.825 0.64 ;
        RECT 1.545 -0.18 1.785 0.32 ;
        RECT 0.135 -0.18 0.255 0.885 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.54 2.79 ;
        RECT 6.57 1.98 6.69 2.79 ;
        RECT 4.06 2.22 4.3 2.79 ;
        RECT 3.52 2.16 3.64 2.79 ;
        RECT 1.425 2.04 1.545 2.79 ;
        RECT 0.135 1.845 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.935 1.345 6.85 1.345 6.85 1.86 5.83 1.86 5.83 2.03 5.59 2.03 5.59 1.86 5.38 1.86 5.38 2 5.26 2 5.26 1.74 6.73 1.74 6.73 0.88 6.515 0.88 6.515 0.58 5.445 0.58 5.445 0.46 6.635 0.46 6.635 0.76 6.85 0.76 6.85 1.105 6.935 1.105 ;
      POLYGON 5.265 0.58 5.145 0.58 5.145 0.66 4.185 0.66 4.185 0.58 4.065 0.58 4.065 0.46 4.305 0.46 4.305 0.54 5.025 0.54 5.025 0.46 5.265 0.46 ;
      POLYGON 5.16 1.62 5.14 1.62 5.14 2.18 4.42 2.18 4.42 2.1 3.85 2.1 3.85 2.04 3.585 2.04 3.585 2.03 2.79 2.03 2.79 1.96 1.665 1.96 1.665 1.92 0.825 1.92 0.825 1.365 0.515 1.365 0.515 1.485 0.395 1.485 0.395 1.245 0.825 1.245 0.825 0.44 2.385 0.44 2.385 0.41 3.125 0.41 3.125 0.46 3.245 0.46 3.245 0.58 3.005 0.58 3.005 0.53 2.505 0.53 2.505 0.9 2.385 0.9 2.385 0.56 0.945 0.56 0.945 1.8 1.785 1.8 1.785 1.84 2.385 1.84 2.385 1.66 2.505 1.66 2.505 1.84 2.79 1.84 2.79 1.79 2.91 1.79 2.91 1.91 3.705 1.91 3.705 1.92 3.97 1.92 3.97 1.98 4.54 1.98 4.54 2.06 5.02 2.06 5.02 1.62 4.92 1.62 4.92 1.5 5.16 1.5 ;
      POLYGON 4.9 1.94 4.66 1.94 4.66 1.8 3.88 1.8 3.88 1.56 4 1.56 4 1.68 4.78 1.68 4.78 1.82 4.9 1.82 ;
      POLYGON 2.145 0.84 1.245 0.84 1.245 0.92 1.125 0.92 1.125 0.68 1.245 0.68 1.245 0.72 2.145 0.72 ;
      POLYGON 2.145 1.72 1.905 1.72 1.905 1.68 1.065 1.68 1.065 1.56 2.025 1.56 2.025 1.6 2.145 1.6 ;
  END
END ADDFXL

MACRO INVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX6 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.84 1.15 1.4 1.27 ;
        RECT 0.885 1.15 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.32 1.43 2.44 2.21 ;
        RECT 0.58 0.91 2.44 1.03 ;
        RECT 2.32 0.4 2.44 1.03 ;
        RECT 0.64 1.5 2.44 1.62 ;
        RECT 1.52 1.175 1.67 1.62 ;
        RECT 1.52 0.91 1.64 1.62 ;
        RECT 1.48 1.43 1.6 2.21 ;
        RECT 1.48 0.4 1.6 1.03 ;
        RECT 0.64 1.43 0.76 2.21 ;
        RECT 0.58 0.4 0.7 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.9 -0.18 2.02 0.79 ;
        RECT 1.06 -0.18 1.18 0.79 ;
        RECT 0.16 -0.18 0.28 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.9 1.74 2.02 2.79 ;
        RECT 1.06 1.74 1.18 2.79 ;
        RECT 0.22 1.43 0.34 2.79 ;
    END
  END VDD
END INVX6

MACRO AOI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.005 0.935 1.25 ;
        RECT 0.65 1.005 0.935 1.145 ;
        RECT 0.65 0.88 0.8 1.145 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 1 1.38 1.435 ;
        RECT 1.21 1 1.33 1.46 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1 1.67 1.475 ;
        RECT 1.52 1 1.67 1.45 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.97 0.51 1.44 ;
        RECT 0.39 0.94 0.51 1.44 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3196 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.885 1.96 1.145 ;
        RECT 1.815 0.76 1.935 2.21 ;
        RECT 1.81 0.76 1.935 1.145 ;
        RECT 1.295 0.76 1.935 0.88 ;
        RECT 1.295 0.59 1.415 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.715 -0.18 1.835 0.64 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 0.975 1.82 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 2.21 1.395 2.21 1.395 1.715 1.215 1.715 1.215 1.7 0.675 1.7 0.675 2.21 0.555 2.21 0.555 1.56 0.675 1.56 0.675 1.58 1.335 1.58 1.335 1.595 1.515 1.595 ;
  END
END AOI31X1

MACRO NAND3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.785 0.51 1.24 ;
        RECT 0.36 0.76 0.48 1.24 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 0.93 0.935 1.17 ;
        RECT 0.65 0.93 0.935 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1 1.67 1.5 ;
        RECT 1.52 1 1.67 1.47 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5104 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.36 1.095 2.21 ;
        RECT 0.12 1.36 1.095 1.48 ;
        RECT 0.12 0.52 0.455 0.64 ;
        RECT 0.335 0.4 0.455 0.64 ;
        RECT 0.135 1.36 0.255 2.21 ;
        RECT 0.07 1.175 0.24 1.435 ;
        RECT 0.12 0.52 0.24 1.48 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.295 -0.18 1.415 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.395 1.62 1.515 2.79 ;
        RECT 0.555 1.6 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.995 1.8 1.875 1.8 1.875 1.68 1.79 1.68 1.79 0.88 1.4 0.88 1.4 1.11 1.15 1.11 1.15 0.99 1.28 0.99 1.28 0.76 1.775 0.76 1.775 0.59 1.895 0.59 1.895 0.71 1.91 0.71 1.91 1.56 1.995 1.56 ;
  END
END NAND3BX1

MACRO AO21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.205 1.105 1.38 1.435 ;
        RECT 1.195 1 1.34 1.325 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 0.72 0.88 0.96 ;
        RECT 0.65 0.595 0.84 0.855 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.76 0.51 1.26 ;
        RECT 0.36 0.76 0.51 1.23 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.15 1.295 2.27 2.21 ;
        RECT 1.81 1.295 2.27 1.415 ;
        RECT 1.81 1.175 1.96 1.435 ;
        RECT 1.84 0.59 1.96 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.42 -0.18 1.54 0.64 ;
        RECT 0.26 -0.18 0.38 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.73 1.945 1.85 2.79 ;
        RECT 0.58 1.62 0.7 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.68 1.23 1.62 1.23 1.62 1.675 1.54 1.675 1.54 1.795 1.42 1.795 1.42 1.555 1.5 1.555 1.5 0.88 1 0.88 1 0.4 1.12 0.4 1.12 0.76 1.62 0.76 1.62 0.99 1.68 0.99 ;
      POLYGON 1.18 1.68 0.82 1.68 0.82 1.5 0.34 1.5 0.34 1.68 0.1 1.68 0.1 1.56 0.22 1.56 0.22 1.38 0.94 1.38 0.94 1.56 1.18 1.56 ;
  END
END AO21X1

MACRO OAI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.065 2.29 1.435 ;
        RECT 2.17 1.06 2.29 1.435 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.98 1.96 1.435 ;
        RECT 1.81 0.98 1.93 1.465 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 1.365 0.9 1.635 ;
        RECT 0.65 1.465 0.8 1.75 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 1.255 1.435 1.41 ;
        RECT 1.11 1.22 1.435 1.41 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.51 1.595 ;
        RECT 0.36 0.96 0.48 1.595 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.312 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.53 0.68 2.65 0.92 ;
        RECT 2.39 1.755 2.54 2.015 ;
        RECT 2.29 1.585 2.53 1.945 ;
        RECT 2.41 0.8 2.53 2.015 ;
        RECT 1.02 1.585 2.53 1.705 ;
        RECT 1.02 1.585 1.14 1.945 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1 -0.18 1.12 0.53 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.66 1.825 1.78 2.79 ;
        RECT 0.3 1.825 0.42 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.23 0.92 2.11 0.92 2.11 0.62 1.45 0.62 1.45 0.86 1.21 0.86 1.21 0.74 1.33 0.74 1.33 0.5 2.23 0.5 ;
      POLYGON 1.87 0.86 1.69 0.86 1.69 1.1 0.63 1.1 0.63 0.84 0.46 0.84 0.46 0.72 0.75 0.72 0.75 0.98 1.57 0.98 1.57 0.74 1.87 0.74 ;
  END
END OAI221XL

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1 0.8 1.455 ;
        RECT 0.65 1 0.77 1.48 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.885 0.51 1.29 ;
        RECT 0.33 0.91 0.45 1.33 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 1.13 1.11 1.555 ;
        RECT 0.94 1.175 1.09 1.58 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.44 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 0.76 1.515 0.88 ;
        RECT 1.395 0.59 1.515 0.88 ;
        RECT 1.23 1.175 1.38 1.435 ;
        RECT 1.23 0.76 1.35 2.1 ;
        RECT 0.555 0.645 0.855 0.765 ;
        RECT 0.555 0.525 0.675 0.765 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.17 1.45 0.29 2.79 ;
    END
  END VDD
END NOR3X1

MACRO AND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X4 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.97 0.51 1.21 ;
        RECT 0.07 0.97 0.51 1.09 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.33 1.09 1.725 ;
        RECT 0.95 1.24 1.07 1.725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 1.51 1.32 2.51 1.44 ;
        RECT 2.39 0.76 2.51 1.44 ;
        RECT 2.35 1.32 2.47 2.21 ;
        RECT 1.57 0.76 2.51 0.88 ;
        RECT 2.35 0.64 2.47 0.88 ;
        RECT 1.45 0.71 1.69 0.83 ;
        RECT 1.51 1.32 1.63 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.77 -0.18 2.89 0.7 ;
        RECT 1.87 0.52 2.11 0.64 ;
        RECT 1.87 -0.18 1.99 0.64 ;
        RECT 1.09 -0.18 1.21 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.77 1.56 2.89 2.79 ;
        RECT 1.93 1.56 2.05 2.79 ;
        RECT 1.09 1.845 1.21 2.79 ;
        RECT 0.25 1.56 0.37 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.27 1.17 2.03 1.17 2.03 1.12 1.85 1.12 1.85 1.17 1.61 1.17 1.61 1.12 0.79 1.12 0.79 2.21 0.67 2.21 0.67 0.83 0.39 0.83 0.39 0.71 0.79 0.71 0.79 1 2.15 1 2.15 1.05 2.27 1.05 ;
  END
END AND2X4

MACRO XOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.18 2.175 1.345 ;
        RECT 1.755 1.18 2.015 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.795 0.94 3.915 1.18 ;
        RECT 3.015 0.97 3.915 1.09 ;
        RECT 3.495 0.94 3.915 1.09 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 1.74 1.575 2.21 ;
        RECT 1.215 0.7 1.515 0.82 ;
        RECT 1.395 0.58 1.515 0.82 ;
        RECT 1.275 1.74 1.575 1.86 ;
        RECT 1.275 1.32 1.395 1.86 ;
        RECT 0.65 0.84 1.335 0.96 ;
        RECT 1.215 0.7 1.335 0.96 ;
        RECT 0.65 1.32 1.395 1.44 ;
        RECT 0.65 1.175 0.8 1.44 ;
        RECT 0.65 0.73 0.77 1.56 ;
        RECT 0.615 1.44 0.735 2.21 ;
        RECT 0.495 0.73 0.77 0.85 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.535 0.46 3.775 0.58 ;
        RECT 3.535 -0.18 3.655 0.58 ;
        RECT 1.815 -0.18 1.935 0.72 ;
        RECT 0.975 -0.18 1.095 0.72 ;
        RECT 0.135 -0.18 0.255 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.595 1.77 3.715 2.79 ;
        RECT 1.815 2.01 2.055 2.15 ;
        RECT 1.815 2.01 1.935 2.79 ;
        RECT 1.035 1.56 1.155 2.79 ;
        RECT 0.195 1.56 0.315 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.155 1.89 4.135 1.89 4.135 2.01 4.015 2.01 4.015 1.77 4.035 1.77 4.035 0.82 2.895 0.82 2.895 1.29 3.275 1.29 3.275 1.41 2.775 1.41 2.775 1.05 2.655 1.05 2.655 1.17 2.535 1.17 2.535 0.93 2.775 0.93 2.775 0.7 4.015 0.7 4.015 0.4 4.135 0.4 4.135 0.52 4.155 0.52 ;
      POLYGON 3.635 1.41 3.515 1.41 3.515 1.65 2.655 1.65 2.655 2.01 2.535 2.01 2.535 1.65 2.295 1.65 2.295 0.65 2.555 0.65 2.555 0.77 2.415 0.77 2.415 1.53 3.395 1.53 3.395 1.29 3.635 1.29 ;
      POLYGON 3.075 2.25 2.175 2.25 2.175 1.89 1.91 1.89 1.91 1.62 1.515 1.62 1.515 1.2 1.255 1.2 1.255 1.08 1.515 1.08 1.515 0.94 2.055 0.94 2.055 0.41 2.855 0.41 2.855 0.46 2.975 0.46 2.975 0.58 2.735 0.58 2.735 0.53 2.175 0.53 2.175 1.06 1.635 1.06 1.635 1.5 2.03 1.5 2.03 1.77 2.295 1.77 2.295 2.13 2.955 2.13 2.955 1.77 3.075 1.77 ;
  END
END XOR2X4

MACRO SDFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX1 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.72 0.36 5.96 0.48 ;
        RECT 5.12 0.83 5.84 0.95 ;
        RECT 5.72 0.36 5.84 0.95 ;
        RECT 5.12 0.38 5.24 0.95 ;
        RECT 3.745 0.38 5.24 0.5 ;
        RECT 3.745 1.23 4.045 1.38 ;
        RECT 3.065 1.29 3.905 1.41 ;
        RECT 3.745 0.38 3.865 1.41 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.53 0.87 8.65 1.33 ;
        RECT 8.48 0.885 8.65 1.32 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.8 1.125 9.05 1.31 ;
        RECT 8.77 0.885 8.92 1.25 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.145 1.23 10.35 1.47 ;
        RECT 9.87 1.23 10.35 1.38 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.55 0.87 10.67 1.11 ;
        RECT 9.63 0.97 10.67 1.09 ;
        RECT 10.01 0.94 10.425 1.09 ;
        RECT 10.01 0.87 10.13 1.11 ;
        RECT 9.41 1.26 9.75 1.38 ;
        RECT 9.63 0.97 9.75 1.38 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 0.74 0.81 0.86 ;
        RECT 0.65 0.74 0.8 1.145 ;
        RECT 0.65 0.74 0.77 1.42 ;
        RECT 0.63 1.3 0.75 1.99 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.98 0.68 2.1 1.585 ;
        RECT 1.92 1.34 2.04 1.99 ;
        RECT 1.81 1.465 2.04 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.49 -0.18 10.61 0.75 ;
        RECT 8.99 -0.18 9.11 0.75 ;
        RECT 6.8 -0.18 6.92 0.63 ;
        RECT 5.36 0.59 5.6 0.71 ;
        RECT 5.48 -0.18 5.6 0.71 ;
        RECT 2.965 -0.18 3.085 0.89 ;
        RECT 1.5 -0.18 1.62 0.73 ;
        RECT 0.15 -0.18 0.27 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.31 1.88 10.43 2.79 ;
        RECT 9.03 1.88 9.15 2.79 ;
        RECT 6.9 2.11 7.02 2.79 ;
        RECT 5.88 2.29 6.12 2.79 ;
        RECT 3.63 2.03 3.87 2.15 ;
        RECT 3.63 2.03 3.75 2.79 ;
        RECT 2.85 1.97 2.97 2.79 ;
        RECT 1.5 1.34 1.62 2.79 ;
        RECT 0.21 1.34 0.33 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.03 0.75 10.91 0.75 10.91 1.83 10.85 1.83 10.85 2 10.73 2 10.73 1.71 9.87 1.71 9.87 1.62 9.75 1.62 9.75 1.5 9.99 1.5 9.99 1.59 10.79 1.59 10.79 0.63 10.91 0.63 10.91 0.51 11.03 0.51 ;
      POLYGON 9.97 0.75 9.51 0.75 9.51 0.99 9.29 0.99 9.29 1.57 9.63 1.57 9.63 1.83 9.79 1.83 9.79 2.07 9.67 2.07 9.67 1.95 9.51 1.95 9.51 1.69 8.12 1.69 8.12 1.57 8.24 1.57 8.24 0.72 8.12 0.72 8.12 0.6 8.36 0.6 8.36 1.57 9.17 1.57 9.17 0.87 9.39 0.87 9.39 0.63 9.85 0.63 9.85 0.51 9.97 0.51 ;
      POLYGON 8.79 1.99 7.62 1.99 7.62 2.15 7.38 2.15 7.38 1.99 6.595 1.99 6.595 2.17 5.56 2.17 5.56 2.05 6.475 2.05 6.475 1.87 7.88 1.87 7.88 0.36 8.69 0.36 8.69 0.75 8.57 0.75 8.57 0.48 8 0.48 8 1.87 8.79 1.87 ;
      POLYGON 7.76 1.35 7.72 1.35 7.72 1.75 7.6 1.75 7.6 1.35 6.6 1.35 6.6 1.23 7.64 1.23 7.64 0.54 7.76 0.54 ;
      POLYGON 7.52 1.06 7.28 1.06 7.28 0.87 6.56 0.87 6.56 0.5 6.2 0.5 6.2 0.72 6.08 0.72 6.08 1.19 5.64 1.19 5.64 1.69 5.4 1.69 5.4 1.57 5.52 1.57 5.52 1.19 4.645 1.19 4.645 1.03 4.88 1.03 4.88 0.62 5 0.62 5 1.07 5.96 1.07 5.96 0.6 6.08 0.6 6.08 0.38 6.68 0.38 6.68 0.75 7.4 0.75 7.4 0.94 7.52 0.94 ;
      POLYGON 7.16 1.11 6.48 1.11 6.48 1.51 6.54 1.51 6.54 1.75 6.01 1.75 6.01 1.93 5.07 1.93 5.07 1.43 4.405 1.43 4.405 0.71 4.645 0.71 4.645 0.83 4.525 0.83 4.525 1.31 5.19 1.31 5.19 1.81 5.89 1.81 5.89 1.63 6.36 1.63 6.36 1.11 6.32 1.11 6.32 0.62 6.44 0.62 6.44 0.99 7.16 0.99 ;
      POLYGON 4.77 1.85 4.65 1.85 4.65 1.67 2.71 1.67 2.71 1.55 4.165 1.55 4.165 0.83 3.985 0.83 3.985 0.71 4.285 0.71 4.285 1.55 4.77 1.55 ;
      POLYGON 4.41 1.91 3.495 1.91 3.495 2.03 3.21 2.03 3.21 1.91 3.375 1.91 3.375 1.79 4.41 1.79 ;
      POLYGON 3.625 1.17 2.59 1.17 2.59 1.91 2.61 1.91 2.61 2.03 2.37 2.03 2.37 1.91 2.47 1.91 2.47 0.77 2.545 0.77 2.545 0.65 2.535 0.65 2.535 0.56 1.86 0.56 1.86 1.18 1.62 1.18 1.62 1.06 1.74 1.06 1.74 0.44 2.655 0.44 2.655 0.53 2.665 0.53 2.665 0.89 2.59 0.89 2.59 1.05 3.625 1.05 ;
      POLYGON 1.14 1.58 1.02 1.58 1.02 0.62 0.45 0.62 0.45 1.06 0.53 1.06 0.53 1.18 0.29 1.18 0.29 1.06 0.33 1.06 0.33 0.5 1.14 0.5 ;
  END
END SDFFSX1

MACRO AOI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X4 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.48 ;
        RECT 0.375 1.01 0.495 1.51 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.01 0.835 1.39 ;
        RECT 0.65 1.065 0.8 1.435 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.365 0.99 7.825 1.11 ;
        RECT 7.365 0.41 7.485 1.11 ;
        RECT 6.565 0.41 7.485 0.53 ;
        RECT 6.565 0.41 6.685 1.09 ;
        RECT 4.945 0.97 6.685 1.09 ;
        RECT 4.945 0.94 5.205 1.09 ;
        RECT 4.925 0.99 5.165 1.11 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.685 1.26 7.005 1.38 ;
        RECT 5.815 1.23 6.075 1.38 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.585 1.5 7.705 2.01 ;
        RECT 4.945 1.5 7.705 1.62 ;
        RECT 7.125 0.65 7.245 1.62 ;
        RECT 6.905 0.65 7.245 0.77 ;
        RECT 6.745 1.5 6.865 2.01 ;
        RECT 5.905 1.5 6.025 2.01 ;
        RECT 5.16 0.65 5.665 0.77 ;
        RECT 2.85 0.7 5.28 0.82 ;
        RECT 4.945 1.5 5.205 1.67 ;
        RECT 5.065 1.5 5.185 2.01 ;
        RECT 4.945 1.23 5.065 1.67 ;
        RECT 4.685 1.23 5.065 1.35 ;
        RECT 4.685 0.7 4.805 1.35 ;
        RECT 3.745 0.65 3.985 0.82 ;
        RECT 2.465 0.65 2.97 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.605 -0.18 7.725 0.64 ;
        RECT 6.325 -0.18 6.445 0.64 ;
        RECT 4.585 0.46 4.825 0.58 ;
        RECT 4.585 -0.18 4.705 0.58 ;
        RECT 3.105 0.46 3.345 0.58 ;
        RECT 3.105 -0.18 3.225 0.58 ;
        RECT 1.885 -0.18 2.005 0.64 ;
        RECT 0.555 -0.18 0.675 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 4.165 1.71 4.405 2.15 ;
        RECT 4.165 1.71 4.285 2.79 ;
        RECT 3.385 1.71 3.505 2.79 ;
        RECT 2.545 1.71 2.665 2.79 ;
        RECT 1.705 1.71 1.825 2.79 ;
        RECT 0.555 1.63 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.125 2.25 4.645 2.25 4.645 1.59 3.925 1.59 3.925 2.21 3.805 2.21 3.805 1.59 3.085 1.59 3.085 2.21 2.965 2.21 2.965 1.59 2.245 1.59 2.245 2.21 2.125 2.21 2.125 1.59 1.405 1.59 1.405 2.21 1.285 2.21 1.285 1.47 4.765 1.47 4.765 2.13 5.485 2.13 5.485 1.74 5.605 1.74 5.605 2.13 6.325 2.13 6.325 1.74 6.445 1.74 6.445 2.13 7.165 2.13 7.165 1.74 7.285 1.74 7.285 2.13 8.005 2.13 8.005 1.56 8.125 1.56 ;
      POLYGON 4.565 1.35 1.155 1.35 1.155 1.68 1.095 1.68 1.095 1.8 0.975 1.8 0.975 1.56 1.035 1.56 1.035 0.6 1.155 0.6 1.155 1.23 4.565 1.23 ;
      POLYGON 3.825 1.11 2.225 1.11 2.225 0.88 1.43 0.88 1.43 0.48 0.915 0.48 0.915 0.89 0.24 0.89 0.24 1.6 0.255 1.6 0.255 2.21 0.135 2.21 0.135 1.72 0.12 1.72 0.12 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.77 0.795 0.77 0.795 0.36 1.55 0.36 1.55 0.76 2.345 0.76 2.345 0.99 3.825 0.99 ;
  END
END AOI2BB2X4

MACRO NOR4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1 0.51 1.475 ;
        RECT 0.36 1 0.51 1.45 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.165 1.145 1.405 ;
        RECT 0.815 1.07 1.055 1.285 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.21 1.725 1.39 ;
        RECT 1.265 1.21 1.725 1.355 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.25 1.53 ;
        RECT 2.1 1.06 2.22 1.56 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4572 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.59 1.575 0.85 ;
        RECT 0.12 0.76 1.555 0.88 ;
        RECT 1.435 0.73 1.575 0.85 ;
        RECT 0.615 0.59 0.735 0.88 ;
        RECT 0.395 1.595 0.515 2.21 ;
        RECT 0.12 1.595 0.515 1.715 ;
        RECT 0.12 0.76 0.24 1.715 ;
        RECT 0.07 0.885 0.24 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.875 -0.18 1.995 0.64 ;
        RECT 1.035 -0.18 1.155 0.64 ;
        RECT 0.195 -0.18 0.315 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.805 1.56 1.925 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.49 1.8 2.405 1.8 2.405 1.92 2.285 1.92 2.285 1.68 2.37 1.68 2.37 0.94 1.915 0.94 1.915 1.09 1.675 1.09 1.675 0.97 1.795 0.97 1.795 0.82 2.355 0.82 2.355 0.59 2.475 0.59 2.475 0.71 2.49 0.71 ;
  END
END NOR4BX1

MACRO SEDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX1 0 0 ;
  SIZE 14.79 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.87 1.13 6.1 1.44 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.2 0.81 8.32 1.2 ;
        RECT 7.115 0.81 8.32 0.93 ;
        RECT 7.115 0.81 7.235 1.2 ;
        RECT 6.975 0.94 7.235 1.09 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.56 1.05 7.76 1.435 ;
        RECT 7.56 1.05 7.68 1.45 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.21 1.35 10.45 1.505 ;
        RECT 10.22 1.35 10.37 1.725 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.41 1.465 13.56 1.725 ;
        RECT 13.41 1.27 13.53 1.725 ;
        RECT 12.47 1.27 13.53 1.39 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 14.24 1.04 14.36 1.28 ;
        RECT 14.02 1.16 14.36 1.28 ;
        RECT 13.99 1.175 14.14 1.435 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.62 1.175 9.79 1.435 ;
        RECT 9.4 1.49 9.74 1.61 ;
        RECT 9.62 0.68 9.74 1.61 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.79 0.18 ;
        RECT 14.1 -0.18 14.22 0.92 ;
        RECT 12.21 0.55 12.45 0.67 ;
        RECT 12.21 -0.18 12.33 0.67 ;
        RECT 11.67 0.55 11.91 0.67 ;
        RECT 11.67 -0.18 11.79 0.67 ;
        RECT 10.55 0.6 10.79 0.72 ;
        RECT 10.67 -0.18 10.79 0.72 ;
        RECT 9.14 -0.18 9.26 0.73 ;
        RECT 7.28 0.33 7.52 0.45 ;
        RECT 7.28 -0.18 7.4 0.45 ;
        RECT 5.8 -0.18 5.92 0.77 ;
        RECT 3.69 0.61 3.93 0.73 ;
        RECT 3.81 -0.18 3.93 0.73 ;
        RECT 1.99 -0.18 2.11 0.86 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.79 2.79 ;
        RECT 14.16 2 14.28 2.79 ;
        RECT 10.4 2.23 10.64 2.79 ;
        RECT 8.92 1.97 9.16 2.09 ;
        RECT 8.92 1.97 9.04 2.79 ;
        RECT 7.28 2.29 7.52 2.79 ;
        RECT 5.8 2.29 6.04 2.79 ;
        RECT 3.87 1.81 3.99 2.79 ;
        RECT 3.75 1.81 3.99 1.93 ;
        RECT 1.85 1.94 2.09 2.06 ;
        RECT 1.85 1.94 1.97 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.655 1.84 13.86 1.84 13.86 2.05 13.05 2.05 13.05 2.19 12.81 2.19 12.81 2.07 12.93 2.07 12.93 1.93 13.74 1.93 13.74 1.72 14.535 1.72 14.535 0.92 14.52 0.92 14.52 0.68 14.64 0.68 14.64 0.8 14.655 0.8 ;
      POLYGON 13.8 1.6 13.68 1.6 13.68 1.15 11.56 1.15 11.56 1.03 13.68 1.03 13.68 0.68 13.8 0.68 ;
      POLYGON 13.13 1.81 13.01 1.81 13.01 1.63 12.29 1.63 12.29 1.81 12.17 1.81 12.17 1.39 11.32 1.39 11.32 0.91 11.15 0.91 11.15 0.96 10.31 0.96 10.31 0.48 9.635 0.48 9.635 0.56 9.5 0.56 9.5 0.97 9.04 0.97 9.04 1.2 8.92 1.2 8.92 0.85 9.38 0.85 9.38 0.44 9.515 0.44 9.515 0.36 10.43 0.36 10.43 0.84 11.03 0.84 11.03 0.54 11.15 0.54 11.15 0.66 11.44 0.66 11.44 0.79 12.585 0.79 12.585 0.55 13.09 0.55 13.09 0.67 12.705 0.67 12.705 0.91 11.44 0.91 11.44 1.27 12.29 1.27 12.29 1.51 13.13 1.51 ;
      POLYGON 12.77 1.87 12.65 1.87 12.65 2.05 12.14 2.05 12.14 2.11 11.38 2.11 11.38 1.99 11.36 1.99 11.36 1.75 11.48 1.75 11.48 1.87 11.5 1.87 11.5 1.99 12.02 1.99 12.02 1.93 12.53 1.93 12.53 1.75 12.77 1.75 ;
      POLYGON 11.9 1.87 11.78 1.87 11.78 1.63 11.06 1.63 11.06 1.87 10.94 1.87 10.94 1.51 11.9 1.51 ;
      POLYGON 11.26 2.25 11.015 2.25 11.015 2.11 9.69 2.11 9.69 1.85 8.8 1.85 8.8 2.17 4.175 2.17 4.175 1.69 3.63 1.69 3.63 2.11 2.45 2.11 2.45 2.25 2.21 2.25 2.21 2.13 2.225 2.13 2.225 1.82 1.55 1.82 1.55 1.87 1.43 1.87 1.43 1.82 1.075 1.82 1.075 1.96 0.835 1.96 0.835 1.84 0.955 1.84 0.955 1.7 1.43 1.7 1.43 1.63 1.57 1.63 1.57 0.62 1.69 0.62 1.69 1.7 2.345 1.7 2.345 1.99 3.51 1.99 3.51 1.57 4.295 1.57 4.295 2.05 8.68 2.05 8.68 1.73 9.16 1.73 9.16 1.21 9.24 1.21 9.24 1.09 9.36 1.09 9.36 1.33 9.28 1.33 9.28 1.73 9.81 1.73 9.81 1.99 11.135 1.99 11.135 2.13 11.26 2.13 ;
      POLYGON 10.84 1.23 10.09 1.23 10.09 1.625 10.1 1.625 10.1 1.87 9.98 1.87 9.98 1.745 9.97 1.745 9.97 0.72 9.95 0.72 9.95 0.6 10.19 0.6 10.19 0.72 10.09 0.72 10.09 1.11 10.84 1.11 ;
      POLYGON 8.76 0.48 7.76 0.48 7.76 0.69 6.855 0.69 6.855 1.57 7.88 1.57 7.88 1.17 8 1.17 8 1.69 6.735 1.69 6.735 0.57 7.64 0.57 7.64 0.36 8.76 0.36 ;
      POLYGON 8.56 1.69 8.24 1.69 8.24 1.93 4.99 1.93 4.99 0.86 4.93 0.86 4.93 0.62 5.05 0.62 5.05 0.74 5.11 0.74 5.11 1.81 8.12 1.81 8.12 1.57 8.44 1.57 8.44 0.62 8.56 0.62 ;
      POLYGON 6.46 1.69 6.34 1.69 6.34 1.57 6.22 1.57 6.22 1.01 5.75 1.01 5.75 1.14 5.63 1.14 5.63 0.89 6.22 0.89 6.22 0.53 6.34 0.53 6.34 1.45 6.46 1.45 ;
      POLYGON 5.5 1.69 5.38 1.69 5.38 0.53 5.17 0.53 5.17 0.5 4.81 0.5 4.81 1.31 4.87 1.31 4.87 1.55 4.75 1.55 4.75 1.43 4.69 1.43 4.69 0.5 4.17 0.5 4.17 0.97 3.45 0.97 3.45 0.5 2.61 0.5 2.61 1.22 2.67 1.22 2.67 1.34 2.43 1.34 2.43 1.22 2.49 1.22 2.49 0.38 3.01 0.38 3.01 0.36 3.25 0.36 3.25 0.38 3.57 0.38 3.57 0.85 4.05 0.85 4.05 0.38 4.25 0.38 4.25 0.36 4.49 0.36 4.49 0.38 5.29 0.38 5.29 0.41 5.5 0.41 ;
      POLYGON 4.57 1.87 4.45 1.87 4.45 1.21 3.47 1.21 3.47 1.09 4.45 1.09 4.45 0.62 4.57 0.62 ;
      POLYGON 4.15 1.45 3.33 1.45 3.33 1.87 3.21 1.87 3.21 0.62 3.33 0.62 3.33 1.33 4.15 1.33 ;
      POLYGON 2.97 0.8 2.91 0.8 2.91 1.87 2.79 1.87 2.79 1.58 1.85 1.58 1.85 1.31 1.97 1.31 1.97 1.46 2.79 1.46 2.79 0.8 2.73 0.8 2.73 0.68 2.97 0.68 ;
      POLYGON 1.155 1.58 1.035 1.58 1.035 1.18 0.375 1.18 0.375 1.06 1.035 1.06 1.035 0.68 1.155 0.68 ;
  END
END SEDFFTRX1

MACRO SEDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX4 0 0 ;
  SIZE 17.4 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.39 1.98 1.41 ;
        RECT 0.9 0.39 1.98 0.51 ;
        RECT 0.3 0.97 1.22 1.09 ;
        RECT 0.9 0.39 1.02 1.09 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.23 0.88 1.47 ;
        RECT 0.595 1.21 0.855 1.47 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.17 1.175 8.34 1.435 ;
        RECT 7.91 1.3 8.34 1.42 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.065 1.47 13.325 1.74 ;
        RECT 13.085 1.34 13.325 1.74 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.275 1.32 16.24 1.44 ;
        RECT 16.12 1.06 16.24 1.44 ;
        RECT 16.02 1.175 16.24 1.44 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.865 1 16.985 1.24 ;
        RECT 16.6 1 16.985 1.145 ;
        RECT 16.6 0.885 16.75 1.145 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.82 0.72 10.02 0.84 ;
        RECT 9.495 1.52 9.615 1.8 ;
        RECT 9.005 1.52 9.615 1.64 ;
        RECT 8.475 1.62 9.265 1.67 ;
        RECT 8.475 1.62 9.16 1.74 ;
        RECT 9.04 0.72 9.16 1.74 ;
        RECT 8.475 1.62 8.715 1.8 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.74 0.72 11.94 0.84 ;
        RECT 11.355 1.62 11.595 1.74 ;
        RECT 10.745 1.52 11.475 1.64 ;
        RECT 10.395 1.62 11.005 1.67 ;
        RECT 10.395 1.62 10.98 1.74 ;
        RECT 10.86 0.72 10.98 1.74 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 17.4 0.18 ;
        RECT 16.685 -0.18 16.805 0.4 ;
        RECT 15.115 0.6 15.355 0.72 ;
        RECT 15.115 -0.18 15.235 0.72 ;
        RECT 14.785 -0.18 14.905 0.4 ;
        RECT 13.59 -0.18 13.83 0.38 ;
        RECT 12.18 -0.18 12.42 0.36 ;
        RECT 11.22 -0.18 11.46 0.36 ;
        RECT 10.26 -0.18 10.5 0.36 ;
        RECT 9.3 -0.18 9.54 0.36 ;
        RECT 8.34 -0.18 8.58 0.36 ;
        RECT 6.985 0.58 7.225 0.7 ;
        RECT 6.985 -0.18 7.105 0.7 ;
        RECT 6.145 0.58 6.385 0.7 ;
        RECT 6.145 -0.18 6.265 0.7 ;
        RECT 4.265 -0.18 4.505 0.32 ;
        RECT 2.14 -0.18 2.26 0.81 ;
        RECT 0.56 -0.18 0.68 0.81 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 17.4 2.79 ;
        RECT 16.605 2.08 16.845 2.2 ;
        RECT 16.605 2.08 16.725 2.79 ;
        RECT 13.265 2.14 13.385 2.79 ;
        RECT 11.835 2.16 12.075 2.28 ;
        RECT 11.835 2.16 11.955 2.79 ;
        RECT 10.875 2.1 11.115 2.22 ;
        RECT 10.875 2.1 10.995 2.79 ;
        RECT 9.915 2.16 10.155 2.28 ;
        RECT 9.915 2.16 10.035 2.79 ;
        RECT 8.955 2.16 9.195 2.28 ;
        RECT 8.955 2.16 9.075 2.79 ;
        RECT 7.995 2.16 8.235 2.28 ;
        RECT 7.995 2.16 8.115 2.79 ;
        RECT 7.125 2.2 7.365 2.79 ;
        RECT 6.185 2.28 6.425 2.79 ;
        RECT 4.025 2.22 4.145 2.79 ;
        RECT 2.34 2.29 2.58 2.79 ;
        RECT 0.62 1.83 0.86 1.95 ;
        RECT 0.62 1.83 0.74 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 17.265 1.86 16.735 1.86 16.735 1.96 16.47 1.96 16.47 2.24 15.615 2.24 15.615 2.12 16.35 2.12 16.35 1.84 16.615 1.84 16.615 1.74 17.145 1.74 17.145 0.68 17.265 0.68 ;
      POLYGON 16.48 1.68 16.145 1.68 16.145 1.56 16.36 1.56 16.36 0.92 16.205 0.92 16.205 0.48 15.605 0.48 15.605 0.96 14.81 0.96 14.81 1.18 14.57 1.18 14.57 1.06 14.69 1.06 14.69 0.84 15.485 0.84 15.485 0.36 16.325 0.36 16.325 0.8 16.48 0.8 ;
      POLYGON 15.995 0.72 15.845 0.72 15.845 1.2 15.155 1.2 15.155 1.56 15.935 1.56 15.935 1.86 15.815 1.86 15.815 1.68 15.155 1.68 15.155 1.8 14.915 1.8 14.915 1.68 15.035 1.68 15.035 1.42 13.565 1.42 13.565 1.98 13.485 1.98 13.485 2.02 12.955 2.02 12.955 2.04 12.04 2.04 12.04 1.98 10.305 1.98 10.305 2.04 7.655 2.04 7.655 2.08 6.065 2.08 6.065 2.24 4.265 2.24 4.265 2.1 3.905 2.1 3.905 2.17 2.14 2.17 2.14 2.15 2.02 2.15 2.02 2.03 2.26 2.03 2.26 2.05 3.785 2.05 3.785 1.98 4.385 1.98 4.385 2.12 5.945 2.12 5.945 1.96 7.535 1.96 7.535 1.92 10.185 1.92 10.185 1.86 12.16 1.86 12.16 1.92 12.835 1.92 12.835 1.9 13.365 1.9 13.365 1.86 13.445 1.86 13.445 1.3 14.19 1.3 14.19 0.86 14.07 0.86 14.07 0.74 14.31 0.74 14.31 1.3 15.035 1.3 15.035 1.08 15.725 1.08 15.725 0.6 15.995 0.6 ;
      POLYGON 15.575 1.92 15.455 1.92 15.455 2.08 14.225 2.08 14.225 1.9 14.105 1.9 14.105 1.78 14.345 1.78 14.345 1.96 15.335 1.96 15.335 1.8 15.575 1.8 ;
      POLYGON 14.705 1.84 14.585 1.84 14.585 1.66 13.985 1.66 13.985 1.78 13.685 1.78 13.685 1.66 13.865 1.66 13.865 1.54 14.705 1.54 ;
      POLYGON 14.45 0.54 14.07 0.54 14.07 0.62 13.35 0.62 13.35 0.56 12.94 0.56 12.94 0.6 12.41 0.6 12.41 1.24 12.29 1.24 12.29 0.6 8.7 0.6 8.7 0.98 8.92 0.98 8.92 1.22 8.58 1.22 8.58 1.46 8.46 1.46 8.46 1.1 8.58 1.1 8.58 0.6 7.54 0.6 7.54 0.94 6.745 0.94 6.745 1.3 6.765 1.3 6.765 1.48 6.885 1.48 6.885 1.6 6.645 1.6 6.645 1.42 6.005 1.42 6.005 1.18 6.125 1.18 6.125 1.3 6.625 1.3 6.625 0.62 6.745 0.62 6.745 0.82 7.42 0.82 7.42 0.48 12.82 0.48 12.82 0.44 13.47 0.44 13.47 0.5 13.95 0.5 13.95 0.42 14.45 0.42 ;
      POLYGON 13.79 1.18 12.945 1.18 12.945 1.78 12.705 1.78 12.705 1.66 12.825 1.66 12.825 0.96 13.11 0.96 13.11 0.68 13.23 0.68 13.23 1.06 13.79 1.06 ;
      POLYGON 12.9 0.84 12.705 0.84 12.705 1.48 12.495 1.48 12.495 1.8 12.375 1.8 12.375 1.48 11.62 1.48 11.62 1.24 11.74 1.24 11.74 1.36 12.585 1.36 12.585 0.72 12.9 0.72 ;
      POLYGON 8.05 1.18 7.79 1.18 7.79 1.68 7.695 1.68 7.695 1.8 7.15 1.8 7.15 1.84 5.825 1.84 5.825 2 4.505 2 4.505 1.68 3.845 1.68 3.845 1.5 3.78 1.5 3.78 1.26 3.9 1.26 3.9 1.38 3.965 1.38 3.965 1.56 4.625 1.56 4.625 1.88 5.105 1.88 5.105 1.44 4.985 1.44 4.985 1.32 5.225 1.32 5.225 1.88 5.705 1.88 5.705 1.18 5.585 1.18 5.585 1.06 5.825 1.06 5.825 1.72 7.03 1.72 7.03 1.68 7.575 1.68 7.575 1.56 7.67 1.56 7.67 1.06 7.81 1.06 7.81 0.72 8.05 0.72 ;
      POLYGON 6.505 1.18 6.385 1.18 6.385 0.94 5.465 0.94 5.465 1.64 5.585 1.64 5.585 1.76 5.345 1.76 5.345 0.62 5.465 0.62 5.465 0.82 6.505 0.82 ;
      POLYGON 5.225 1.12 4.985 1.12 4.985 1 5.105 1 5.105 0.56 4.025 0.56 4.025 0.5 3.42 0.5 3.42 1.5 3.3 1.5 3.3 0.5 2.89 0.5 2.89 0.57 2.68 0.57 2.68 0.69 2.75 0.69 2.75 1.57 2.94 1.57 2.94 1.69 2.63 1.69 2.63 0.81 2.56 0.81 2.56 0.45 2.77 0.45 2.77 0.38 3.705 0.38 3.705 0.36 3.945 0.36 3.945 0.38 4.145 0.38 4.145 0.44 5.225 0.44 ;
      POLYGON 4.985 0.8 4.865 0.8 4.865 1.64 4.985 1.64 4.985 1.76 4.745 1.76 4.745 1.44 4.085 1.44 4.085 1.32 4.745 1.32 4.745 0.68 4.985 0.68 ;
      POLYGON 4.625 1.12 3.66 1.12 3.66 1.62 3.725 1.62 3.725 1.86 3.605 1.86 3.605 1.74 3.54 1.74 3.54 0.68 3.78 0.68 3.78 0.8 3.66 0.8 3.66 1 4.625 1 ;
      POLYGON 3.305 1.93 2.39 1.93 2.39 1.91 1.6 1.91 1.6 1.55 1.62 1.55 1.62 0.75 1.14 0.75 1.14 0.63 1.74 0.63 1.74 1.67 1.72 1.67 1.72 1.79 2.51 1.79 2.51 1.81 3.06 1.81 3.06 0.62 3.18 0.62 3.18 1.62 3.305 1.62 ;
      POLYGON 1.5 1.43 1.48 1.43 1.48 1.71 0.32 1.71 0.32 1.83 0.2 1.83 0.2 1.71 0.06 1.71 0.06 0.69 0.14 0.69 0.14 0.57 0.26 0.57 0.26 0.81 0.18 0.81 0.18 1.59 1.36 1.59 1.36 1.31 1.38 1.31 1.38 1.19 1.5 1.19 ;
  END
END SEDFFTRX4

MACRO OR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.92 2.015 1.12 ;
        RECT 1.755 0.89 1.875 1.24 ;
    END
  END A
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.31 1.175 0.53 1.435 ;
        RECT 0.335 1.06 0.53 1.435 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.035 0.82 1.44 ;
        RECT 0.7 1.02 0.82 1.44 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.08 1.375 1.32 ;
        RECT 0.94 1.175 1.375 1.295 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.175 2.54 1.435 ;
        RECT 2.415 0.68 2.535 1.435 ;
        RECT 2.335 1.295 2.455 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.835 -0.18 2.955 0.73 ;
        RECT 1.995 -0.18 2.115 0.73 ;
        RECT 1.035 -0.18 1.155 0.38 ;
        RECT 0.135 -0.18 0.255 0.9 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.755 1.56 2.875 2.79 ;
        RECT 1.915 1.6 2.035 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.215 1.48 1.635 1.48 1.635 1.68 0.34 1.68 0.34 1.8 0.22 1.8 0.22 1.56 1.515 1.56 1.515 0.9 0.555 0.9 0.555 0.66 0.675 0.66 0.675 0.78 1.515 0.78 1.515 0.66 1.635 0.66 1.635 1.36 2.095 1.36 2.095 1.24 2.215 1.24 ;
  END
END OR4X2

MACRO DFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX2 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 0.925 0.435 1.165 ;
        RECT 0.07 0.885 0.33 1.145 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 1.315 1.545 1.555 ;
        RECT 1.23 1.315 1.545 1.435 ;
        RECT 1.23 1.175 1.38 1.435 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.065 0.68 5.185 1.66 ;
        RECT 4.965 1.54 5.085 2.19 ;
        RECT 5 1.175 5.185 1.66 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.545 -0.18 5.665 0.76 ;
        RECT 4.585 -0.18 4.705 0.73 ;
        RECT 2.845 -0.18 2.965 0.89 ;
        RECT 1.485 -0.18 1.605 0.38 ;
        RECT 0.135 -0.18 0.255 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.385 1.54 5.505 2.79 ;
        RECT 4.545 1.83 4.665 2.79 ;
        RECT 2.785 2.18 3.025 2.3 ;
        RECT 2.785 2.18 2.905 2.79 ;
        RECT 1.265 1.95 1.385 2.79 ;
        RECT 0.135 1.46 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.105 1.42 5.925 1.42 5.925 2.06 5.805 2.06 5.805 1.42 5.305 1.42 5.305 1.18 5.425 1.18 5.425 1.3 5.985 1.3 5.985 0.62 6.105 0.62 ;
      POLYGON 5.865 1.18 5.745 1.18 5.745 1 5.305 1 5.305 0.56 4.945 0.56 4.945 0.97 3.925 0.97 3.925 1.89 4.045 1.89 4.045 2.01 3.805 2.01 3.805 0.72 4.065 0.72 4.065 0.85 4.825 0.85 4.825 0.44 5.425 0.44 5.425 0.88 5.865 0.88 ;
      POLYGON 4.285 2.25 3.145 2.25 3.145 2.06 2.66 2.06 2.66 2.25 1.745 2.25 1.745 1.795 1.11 1.795 1.11 1.915 0.965 1.915 0.965 2.09 0.845 2.09 0.845 1.795 0.99 1.795 0.99 0.84 0.885 0.84 0.885 0.72 1.125 0.72 1.125 0.84 1.11 0.84 1.11 1.675 1.745 1.675 1.745 1.49 1.865 1.49 1.865 2.13 2.54 2.13 2.54 1.94 3.265 1.94 3.265 2.13 4.165 2.13 4.165 1.75 4.045 1.75 4.045 1.51 4.165 1.51 4.165 1.63 4.285 1.63 ;
      POLYGON 4.225 0.5 3.735 0.5 3.735 0.54 3.685 0.54 3.685 1.58 3.565 1.58 3.565 0.54 3.205 0.54 3.205 1.13 2.465 1.13 2.465 1.58 2.225 1.58 2.225 1.46 2.345 1.46 2.345 1.01 2.445 1.01 2.445 0.6 1.845 0.6 1.845 0.62 1.245 0.62 1.245 0.6 0.675 0.6 0.675 1.58 0.555 1.58 0.555 0.48 1.065 0.48 1.065 0.38 1.365 0.38 1.365 0.5 1.725 0.5 1.725 0.48 1.925 0.48 1.925 0.38 2.165 0.38 2.165 0.48 2.565 0.48 2.565 1.01 3.085 1.01 3.085 0.42 3.615 0.42 3.615 0.38 4.225 0.38 ;
      POLYGON 3.625 2.01 3.385 2.01 3.385 1.82 3.325 1.82 3.325 1.37 2.585 1.37 2.585 1.25 3.325 1.25 3.325 0.66 3.445 0.66 3.445 1.7 3.505 1.7 3.505 1.89 3.625 1.89 ;
      POLYGON 3.185 1.82 2.325 1.82 2.325 2.01 1.985 2.01 1.985 0.72 2.325 0.72 2.325 0.84 2.105 0.84 2.105 1.7 3.065 1.7 3.065 1.49 3.185 1.49 ;
  END
END DFFQX2

MACRO AND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X6 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.295 0.75 2.415 1.22 ;
        RECT 0.39 0.75 2.415 0.87 ;
        RECT 0.495 0.75 0.615 1.22 ;
        RECT 0.36 0.885 0.615 1.145 ;
        RECT 0.39 0.75 0.615 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.99 2.095 1.23 ;
        RECT 1.81 0.99 1.96 1.435 ;
        RECT 0.935 0.99 2.095 1.11 ;
        RECT 0.755 1.04 1.055 1.16 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.25 1.555 1.5 ;
        RECT 1.175 1.23 1.435 1.5 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.755 1.39 4.875 2.21 ;
        RECT 4.735 0.4 4.855 0.915 ;
        RECT 3.075 1.39 4.875 1.51 ;
        RECT 4.555 0.795 4.855 0.915 ;
        RECT 2.995 0.91 4.675 1.03 ;
        RECT 3.955 1.175 4.28 1.51 ;
        RECT 3.955 0.91 4.075 1.51 ;
        RECT 3.915 1.39 4.035 2.21 ;
        RECT 3.895 0.4 4.015 1.03 ;
        RECT 3.075 1.39 3.195 2.21 ;
        RECT 2.995 0.4 3.115 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 4.315 -0.18 4.435 0.79 ;
        RECT 3.475 -0.18 3.595 0.79 ;
        RECT 2.455 -0.18 2.695 0.39 ;
        RECT 0.275 0.51 0.515 0.63 ;
        RECT 0.275 -0.18 0.395 0.63 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.335 1.63 4.455 2.79 ;
        RECT 3.495 1.63 3.615 2.79 ;
        RECT 2.655 1.86 2.775 2.79 ;
        RECT 1.815 1.86 1.935 2.79 ;
        RECT 0.975 1.86 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.835 1.27 2.655 1.27 2.655 1.74 2.355 1.74 2.355 2.21 2.235 2.21 2.235 1.74 1.515 1.74 1.515 2.21 1.395 2.21 1.395 1.74 0.675 1.74 0.675 2.21 0.555 2.21 0.555 1.56 0.675 1.56 0.675 1.62 2.235 1.62 2.235 1.56 2.355 1.56 2.355 1.62 2.535 1.62 2.535 0.63 1.435 0.63 1.435 0.51 2.655 0.51 2.655 1.15 3.835 1.15 ;
  END
END AND3X6

MACRO AOI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X4 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.695 0.99 8.495 1.11 ;
        RECT 7.695 0.94 7.815 1.18 ;
        RECT 7.555 0.94 7.815 1.09 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.155 0.99 7.135 1.11 ;
        RECT 6.685 1.23 6.945 1.38 ;
        RECT 6.685 0.99 6.805 1.38 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.505 0.99 3.505 1.11 ;
        RECT 0.885 0.94 1.145 1.11 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.995 1.23 6.395 1.35 ;
        RECT 5.815 1.23 6.075 1.38 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.345 1.23 2.865 1.35 ;
        RECT 1.465 1.23 1.725 1.38 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2416 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.575 1.32 8.695 2.01 ;
        RECT 7.735 1.32 8.695 1.44 ;
        RECT 8.215 0.65 8.455 0.77 ;
        RECT 1.625 0.7 8.335 0.82 ;
        RECT 7.735 1.32 7.855 2.01 ;
        RECT 3.915 1.5 7.855 1.62 ;
        RECT 7.375 0.65 7.615 0.82 ;
        RECT 6.315 0.65 6.555 0.82 ;
        RECT 4.735 0.65 4.975 0.82 ;
        RECT 3.785 1.23 4.045 1.38 ;
        RECT 3.915 0.7 4.035 1.62 ;
        RECT 2.785 0.65 3.025 0.82 ;
        RECT 1.505 0.65 1.745 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 8.695 -0.18 8.815 0.64 ;
        RECT 7.795 0.46 8.035 0.58 ;
        RECT 7.795 -0.18 7.915 0.58 ;
        RECT 6.955 0.46 7.195 0.58 ;
        RECT 6.955 -0.18 7.075 0.58 ;
        RECT 5.475 0.46 5.715 0.58 ;
        RECT 5.475 -0.18 5.595 0.58 ;
        RECT 3.895 0.46 4.135 0.58 ;
        RECT 3.895 -0.18 4.015 0.58 ;
        RECT 2.145 0.46 2.385 0.58 ;
        RECT 2.145 -0.18 2.265 0.58 ;
        RECT 0.925 -0.18 1.045 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 3.505 1.98 3.745 2.15 ;
        RECT 3.505 1.98 3.625 2.79 ;
        RECT 2.665 1.98 2.905 2.15 ;
        RECT 2.665 1.98 2.785 2.79 ;
        RECT 1.825 1.98 2.065 2.15 ;
        RECT 1.825 1.98 1.945 2.79 ;
        RECT 0.985 1.98 1.225 2.15 ;
        RECT 0.985 1.98 1.105 2.79 ;
        RECT 0.205 1.56 0.325 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.115 2.25 4.015 2.25 4.015 2.15 3.895 2.15 3.895 1.98 4.135 1.98 4.135 2.13 4.735 2.13 4.735 1.98 4.975 1.98 4.975 2.13 5.575 2.13 5.575 1.98 5.815 1.98 5.815 2.13 6.415 2.13 6.415 1.98 6.655 1.98 6.655 2.13 7.315 2.13 7.315 1.74 7.435 1.74 7.435 2.13 8.155 2.13 8.155 1.56 8.275 1.56 8.275 2.13 8.995 2.13 8.995 1.56 9.115 1.56 ;
      POLYGON 7.015 2.01 6.895 2.01 6.895 1.86 6.175 1.86 6.175 2.01 6.055 2.01 6.055 1.86 5.335 1.86 5.335 2.01 5.215 2.01 5.215 1.86 4.495 1.86 4.495 2.01 4.375 2.01 4.375 1.86 3.265 1.86 3.265 2.21 3.145 2.21 3.145 1.86 2.425 1.86 2.425 2.21 2.305 2.21 2.305 1.86 1.585 1.86 1.585 2.21 1.465 2.21 1.465 1.86 0.745 1.86 0.745 2.21 0.625 2.21 0.625 1.56 0.745 1.56 0.745 1.74 1.465 1.74 1.465 1.56 1.585 1.56 1.585 1.74 2.305 1.74 2.305 1.56 2.425 1.56 2.425 1.74 3.145 1.74 3.145 1.56 3.265 1.56 3.265 1.74 7.015 1.74 ;
  END
END AOI221X4

MACRO XOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X2 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 1.22 1.335 1.46 ;
        RECT 0.885 1.23 1.335 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.18 3.175 1.3 ;
        RECT 2.335 1.18 2.595 1.38 ;
        RECT 2.255 1.14 2.495 1.3 ;
        RECT 1.695 1.34 1.935 1.46 ;
        RECT 1.815 1.18 1.935 1.46 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.74 0.715 2.21 ;
        RECT 0.405 0.74 0.675 0.86 ;
        RECT 0.555 0.62 0.675 0.86 ;
        RECT 0.405 1.74 0.715 1.86 ;
        RECT 0.405 0.74 0.525 1.86 ;
        RECT 0.36 0.885 0.525 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.735 -0.18 2.855 0.78 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.615 1.74 2.735 2.79 ;
        RECT 1.015 2.22 1.255 2.79 ;
        RECT 0.165 1.56 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.415 1.74 3.155 1.74 3.155 1.86 3.035 1.86 3.035 1.62 2.335 1.62 2.335 2.24 2.055 2.24 2.055 2.12 2.215 2.12 2.215 1.5 3.155 1.5 3.155 1.62 3.295 1.62 3.295 0.78 3.155 0.78 3.155 0.54 3.275 0.54 3.275 0.66 3.415 0.66 ;
      POLYGON 2.855 1.06 2.615 1.06 2.615 1.02 1.575 1.02 1.575 1.58 1.675 1.58 1.675 1.86 1.555 1.86 1.555 1.7 1.455 1.7 1.455 0.6 1.695 0.6 1.695 0.72 1.575 0.72 1.575 0.9 2.735 0.9 2.735 0.94 2.855 0.94 ;
      POLYGON 2.215 0.78 2.095 0.78 2.095 0.48 1.335 0.48 1.335 1.1 0.765 1.1 0.765 1.5 0.955 1.5 0.955 1.58 1.14 1.58 1.14 1.98 1.815 1.98 1.815 1.86 1.975 1.86 1.975 1.74 2.095 1.74 2.095 1.98 1.935 1.98 1.935 2.1 1.02 2.1 1.02 1.7 0.835 1.7 0.835 1.62 0.645 1.62 0.645 0.98 1.215 0.98 1.215 0.36 2.215 0.36 ;
  END
END XOR2X2

MACRO TLATNCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX12 0 0 ;
  SIZE 10.73 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.23 0.855 1.38 ;
        RECT 0.595 1.08 0.715 1.38 ;
        RECT 0.355 1.08 0.715 1.2 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.93 1.465 10.08 1.725 ;
        RECT 9.93 1.34 10.05 1.725 ;
        RECT 9.895 1.22 10.015 1.46 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.275 1.4 4.515 1.58 ;
        RECT 1.215 0.84 4.515 0.96 ;
        RECT 4.395 0.4 4.515 0.96 ;
        RECT 1.215 1.32 4.395 1.44 ;
        RECT 3.435 1.32 3.675 1.58 ;
        RECT 3.555 0.4 3.675 0.96 ;
        RECT 2.595 1.32 2.835 1.58 ;
        RECT 2.715 0.4 2.835 0.96 ;
        RECT 1.755 1.32 1.995 1.58 ;
        RECT 1.875 0.4 1.995 0.96 ;
        RECT 1.215 1.175 1.38 1.44 ;
        RECT 0.975 1.34 1.335 1.46 ;
        RECT 1.215 0.8 1.335 1.46 ;
        RECT 1.035 0.8 1.335 0.92 ;
        RECT 1.035 0.4 1.155 0.92 ;
        RECT 0.975 1.34 1.095 1.58 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.73 0.18 ;
        RECT 9.975 0.5 10.215 0.62 ;
        RECT 10.095 -0.18 10.215 0.62 ;
        RECT 8.075 -0.18 8.195 0.73 ;
        RECT 6.415 0.55 6.655 0.67 ;
        RECT 6.415 -0.18 6.535 0.67 ;
        RECT 4.815 -0.18 4.935 0.915 ;
        RECT 3.975 -0.18 4.095 0.72 ;
        RECT 3.135 -0.18 3.255 0.72 ;
        RECT 2.295 -0.18 2.415 0.72 ;
        RECT 1.455 -0.18 1.575 0.72 ;
        RECT 0.615 -0.18 0.735 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.73 2.79 ;
        RECT 10.055 1.845 10.175 2.79 ;
        RECT 8.335 2.2 8.455 2.79 ;
        RECT 7.315 2.1 7.555 2.22 ;
        RECT 7.315 2.1 7.435 2.79 ;
        RECT 6.355 2.1 6.595 2.22 ;
        RECT 6.355 2.1 6.475 2.79 ;
        RECT 5.395 2.12 5.635 2.24 ;
        RECT 5.395 2.12 5.515 2.79 ;
        RECT 4.755 2.12 4.995 2.24 ;
        RECT 4.755 2.12 4.875 2.79 ;
        RECT 3.855 1.94 4.095 2.06 ;
        RECT 3.855 1.94 3.975 2.79 ;
        RECT 3.015 1.94 3.255 2.06 ;
        RECT 3.015 1.94 3.135 2.79 ;
        RECT 2.175 1.94 2.415 2.06 ;
        RECT 2.175 1.94 2.295 2.79 ;
        RECT 1.335 1.94 1.575 2.06 ;
        RECT 1.335 1.94 1.455 2.79 ;
        RECT 0.495 1.98 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.595 2.21 10.475 2.21 10.475 1.68 10.455 1.68 10.455 0.86 9.735 0.86 9.735 0.57 8.435 0.57 8.435 1.16 8.315 1.16 8.315 1.18 8.075 1.18 8.075 1.16 6.915 1.16 6.915 1.2 6.675 1.2 6.675 1.04 8.315 1.04 8.315 0.45 9.855 0.45 9.855 0.74 10.455 0.74 10.455 0.63 10.575 0.63 10.575 1.56 10.595 1.56 ;
      POLYGON 10.335 1.22 10.215 1.22 10.215 1.1 9.775 1.1 9.775 1.7 9.535 1.7 9.535 1.74 9.295 1.74 9.295 1.62 9.415 1.62 9.415 1.58 9.655 1.58 9.655 1.1 9.115 1.1 9.115 0.81 8.975 0.81 8.975 0.69 9.235 0.69 9.235 0.98 10.335 0.98 ;
      POLYGON 9.535 1.46 9.415 1.46 9.415 1.44 5.415 1.44 5.415 1.52 5.115 1.52 5.115 1.4 5.295 1.4 5.295 0.675 5.415 0.675 5.415 1.32 5.595 1.32 5.595 1.3 5.835 1.3 5.835 1.32 7.035 1.32 7.035 1.28 7.275 1.28 7.275 1.32 8.875 1.32 8.875 0.97 8.995 0.97 8.995 1.32 9.415 1.32 9.415 1.22 9.535 1.22 ;
      POLYGON 9.195 2.24 9.075 2.24 9.075 2.12 9.03 2.12 9.03 2.08 8.235 2.08 8.235 1.98 6.235 1.98 6.235 2 4.545 2 4.545 1.82 0.135 1.82 0.135 1.58 0.115 1.58 0.115 0.8 0.135 0.8 0.135 0.68 0.255 0.68 0.255 0.92 0.235 0.92 0.235 1.46 0.255 1.46 0.255 1.7 4.665 1.7 4.665 1.88 6.115 1.88 6.115 1.86 8.355 1.86 8.355 1.96 9.15 1.96 9.15 2 9.195 2 ;
      POLYGON 8.035 1.74 5.75 1.74 5.75 1.76 4.875 1.76 4.875 1.2 4.195 1.2 4.195 1.08 5.055 1.08 5.055 0.435 5.705 0.435 5.705 0.55 5.95 0.55 5.95 0.79 6.89 0.79 6.89 0.74 7.395 0.74 7.395 0.86 7.01 0.86 7.01 0.91 5.83 0.91 5.83 0.67 5.585 0.67 5.585 0.555 5.175 0.555 5.175 1.2 4.995 1.2 4.995 1.64 5.63 1.64 5.63 1.62 8.035 1.62 ;
  END
END TLATNCAX12

MACRO AOI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X1 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.76 2.8 2.01 ;
        RECT 2.39 0.76 2.8 0.88 ;
        RECT 2.2 0.65 2.54 0.77 ;
        RECT 2.39 0.595 2.54 0.88 ;
    END
  END Y
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.44 1.025 0.8 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
        RECT 0.44 1.025 0.56 1.265 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.76 1.265 0.88 1.565 ;
        RECT 0.65 1.415 0.8 1.725 ;
    END
  END A0N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.025 2.54 1.48 ;
        RECT 2.42 1 2.54 1.48 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.885 3.12 1.355 ;
        RECT 2.96 0.9 3.08 1.4 ;
    END
  END B0
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.9 -0.18 3.02 0.64 ;
        RECT 1.62 -0.18 1.74 0.64 ;
        RECT 0.66 -0.18 0.78 0.525 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 1.84 1.84 1.96 2.79 ;
        RECT 0.6 1.845 0.72 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.22 2.21 3.175 2.21 3.175 2.25 2.26 2.25 2.26 1.72 1.54 1.72 1.54 2.21 1.42 2.21 1.42 1.56 1.54 1.56 1.54 1.6 2.38 1.6 2.38 2.13 3.055 2.13 3.055 2.09 3.1 2.09 3.1 1.56 3.22 1.56 ;
      POLYGON 2.22 1.17 1.96 1.17 1.96 0.88 1.38 0.88 1.38 0.48 1.02 0.48 1.02 0.765 0.3 0.765 0.3 1.965 0.18 1.965 0.18 0.6 0.3 0.6 0.3 0.645 0.9 0.645 0.9 0.36 1.5 0.36 1.5 0.76 2.08 0.76 2.08 0.93 2.22 0.93 ;
      POLYGON 1.76 1.32 1.26 1.32 1.26 1.845 1.14 1.845 1.14 1.965 1.02 1.965 1.02 1.725 1.14 1.725 1.14 0.6 1.26 0.6 1.26 1.2 1.76 1.2 ;
  END
END AOI2BB2X1

MACRO AND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X8 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.97 2.08 1.09 ;
        RECT 1.84 0.595 1.96 1.09 ;
        RECT 1.81 0.595 1.96 0.855 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.09 ;
        RECT 1.295 1.21 2.78 1.33 ;
        RECT 2.66 0.94 2.78 1.33 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.02 1.105 3.295 1.345 ;
        RECT 0.94 1.45 3.14 1.57 ;
        RECT 3.02 1.105 3.14 1.57 ;
        RECT 0.94 1.175 1.09 1.57 ;
        RECT 0.755 1.28 1.09 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.495 1.69 3.615 1.81 ;
        RECT 3.495 1.22 3.615 1.81 ;
        RECT 3.26 1.465 3.615 1.81 ;
        RECT 0.495 1.22 0.615 1.81 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.915 1.275 7.035 2.21 ;
        RECT 4.395 1.275 7.035 1.395 ;
        RECT 6.595 0.715 6.835 0.835 ;
        RECT 4.135 0.765 6.715 0.885 ;
        RECT 6.075 1.175 6.31 1.435 ;
        RECT 6.075 0.765 6.195 2.21 ;
        RECT 5.755 0.715 5.995 0.885 ;
        RECT 5.235 1.275 5.355 2.21 ;
        RECT 4.915 0.715 5.155 0.885 ;
        RECT 4.395 1.275 4.515 2.21 ;
        RECT 4.015 0.715 4.255 0.835 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.235 -0.18 6.355 0.645 ;
        RECT 5.395 -0.18 5.515 0.645 ;
        RECT 4.495 -0.18 4.615 0.64 ;
        RECT 3.595 0.46 3.835 0.58 ;
        RECT 3.595 -0.18 3.715 0.58 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 6.495 1.515 6.615 2.79 ;
        RECT 5.655 1.515 5.775 2.79 ;
        RECT 4.815 1.515 4.935 2.79 ;
        RECT 3.855 2.17 4.095 2.29 ;
        RECT 3.855 2.17 3.975 2.79 ;
        RECT 2.895 2.17 3.135 2.29 ;
        RECT 2.895 2.17 3.015 2.79 ;
        RECT 1.935 2.17 2.175 2.29 ;
        RECT 1.935 2.17 2.055 2.79 ;
        RECT 0.975 2.17 1.215 2.29 ;
        RECT 0.975 2.17 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.715 1.155 3.855 1.155 3.855 2.05 3.555 2.05 3.555 2.21 3.435 2.21 3.435 2.05 2.595 2.05 2.595 2.21 2.475 2.21 2.475 2.05 1.635 2.05 1.635 2.21 1.515 2.21 1.515 2.05 0.675 2.05 0.675 2.21 0.555 2.21 0.555 1.93 3.735 1.93 3.735 0.82 2.24 0.82 2.24 0.77 2.12 0.77 2.12 0.65 2.36 0.65 2.36 0.7 3.855 0.7 3.855 1.035 5.715 1.035 ;
  END
END AND4X8

MACRO SDFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRXL 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 2.095 1.675 ;
        RECT 1.975 1.32 2.095 1.675 ;
        RECT 1.81 1.465 1.96 1.815 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3012 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.51 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.915 1.25 3.335 1.415 ;
        RECT 2.915 1.23 3.175 1.43 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.035 0.76 8.155 1.03 ;
        RECT 7.9 0.86 8.05 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 0.96 9.575 1.2 ;
        RECT 9.295 0.94 9.555 1.2 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.875 0.94 10.135 1.09 ;
        RECT 9.795 0.7 9.93 1.06 ;
        RECT 8.655 0.7 9.93 0.82 ;
        RECT 9.055 0.7 9.175 0.98 ;
        RECT 8.515 1.1 8.775 1.22 ;
        RECT 8.655 0.7 8.775 1.22 ;
        RECT 8.515 1.1 8.635 1.34 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 1.465 1.67 1.725 ;
        RECT 1.375 0.68 1.495 0.96 ;
        RECT 1.335 0.84 1.455 2.09 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 9.475 0.46 9.715 0.58 ;
        RECT 9.475 -0.18 9.595 0.58 ;
        RECT 8.035 -0.18 8.155 0.64 ;
        RECT 5.355 -0.18 5.595 0.37 ;
        RECT 3.295 0.49 3.535 0.61 ;
        RECT 3.295 -0.18 3.415 0.61 ;
        RECT 1.775 -0.18 1.895 0.4 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 9.535 1.56 9.655 2.79 ;
        RECT 8.095 2.08 8.215 2.79 ;
        RECT 5.995 2.15 6.115 2.79 ;
        RECT 5.095 2.29 5.335 2.79 ;
        RECT 3.465 2.29 3.705 2.79 ;
        RECT 2.565 2.05 2.685 2.79 ;
        RECT 1.755 1.97 1.875 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.375 1.56 10.075 1.56 10.075 1.68 9.955 1.68 9.955 1.44 9.015 1.44 9.015 1.3 8.895 1.3 8.895 1.18 9.135 1.18 9.135 1.32 10.255 1.32 10.255 0.58 9.895 0.58 9.895 0.46 10.375 0.46 ;
      POLYGON 9.075 0.58 8.535 0.58 8.535 0.98 8.395 0.98 8.395 1.5 8.855 1.5 8.855 1.62 8.395 1.62 8.395 1.86 7.225 1.86 7.225 1.36 6.895 1.36 6.895 0.62 7.015 0.62 7.015 1.24 7.345 1.24 7.345 1.74 8.275 1.74 8.275 0.86 8.415 0.86 8.415 0.46 9.075 0.46 ;
      POLYGON 7.955 2.1 6.645 2.1 6.645 2.08 6.38 2.08 6.38 2.03 5.85 2.03 5.85 1.93 2.375 1.93 2.375 1.97 2.295 1.97 2.295 2.09 2.175 2.09 2.175 1.81 2.255 1.81 2.255 0.68 2.375 0.68 2.375 1.81 3.895 1.81 3.895 0.97 4.035 0.97 4.035 1.21 4.015 1.21 4.015 1.81 4.495 1.81 4.495 1.37 4.435 1.37 4.435 1.25 4.675 1.25 4.675 1.37 4.615 1.37 4.615 1.81 5.97 1.81 5.97 1.91 6.5 1.91 6.5 1.96 6.645 1.96 6.645 1.84 6.765 1.84 6.765 1.98 7.955 1.98 ;
      POLYGON 7.795 1.62 7.555 1.62 7.555 1 7.355 1 7.355 1.12 7.235 1.12 7.235 0.5 6.295 0.5 6.295 0.61 5.115 0.61 5.115 0.56 4.635 0.56 4.635 0.97 4.975 0.97 4.975 1.21 4.855 1.21 4.855 1.09 4.515 1.09 4.515 0.44 5.235 0.44 5.235 0.49 6.175 0.49 6.175 0.36 6.415 0.36 6.415 0.38 7.355 0.38 7.355 0.88 7.555 0.88 7.555 0.4 7.675 0.4 7.675 1.5 7.795 1.5 ;
      POLYGON 6.925 1.72 6.805 1.72 6.805 1.6 6.625 1.6 6.625 1.36 5.335 1.36 5.335 0.97 5.455 0.97 5.455 1.24 6.475 1.24 6.475 0.62 6.595 0.62 6.595 1.24 6.745 1.24 6.745 1.48 6.925 1.48 ;
      POLYGON 6.505 1.72 6.385 1.72 6.385 1.69 5.575 1.69 5.575 1.57 6.385 1.57 6.385 1.48 6.505 1.48 ;
      POLYGON 6.155 1.12 5.915 1.12 5.915 0.85 5.215 0.85 5.215 1.69 4.735 1.69 4.735 1.57 5.095 1.57 5.095 0.85 4.755 0.85 4.755 0.68 4.995 0.68 4.995 0.73 6.035 0.73 6.035 1 6.155 1 ;
      RECT 3.145 2.05 5.655 2.17 ;
      POLYGON 4.375 1.69 4.135 1.69 4.135 1.57 4.155 1.57 4.155 0.85 2.895 0.85 2.895 0.48 2.735 0.48 2.735 0.36 3.015 0.36 3.015 0.73 4.155 0.73 4.155 0.62 4.275 0.62 4.275 1.57 4.375 1.57 ;
      POLYGON 3.755 1.14 3.455 1.14 3.455 1.11 2.795 1.11 2.795 1.57 3.225 1.57 3.225 1.69 2.675 1.69 2.675 1.11 2.655 1.11 2.655 0.74 2.495 0.74 2.495 0.56 2.135 0.56 2.135 1.2 1.575 1.2 1.575 1.08 2.015 1.08 2.015 0.44 2.615 0.44 2.615 0.62 2.775 0.62 2.775 0.99 3.575 0.99 3.575 1.02 3.755 1.02 ;
      POLYGON 1.215 1.58 1.095 1.58 1.095 1.46 0.985 1.46 0.985 1.18 0.375 1.18 0.375 1.06 0.985 1.06 0.985 0.68 1.105 0.68 1.105 1.34 1.215 1.34 ;
  END
END SDFFRXL

MACRO XNOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3XL 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 1.35 6.81 1.47 ;
        RECT 6.08 1.23 6.365 1.47 ;
        RECT 6.08 0.905 6.2 1.47 ;
        RECT 5.695 0.905 6.2 1.025 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.252 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.845 0.975 1.025 1.375 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.07 0.325 1.47 ;
        RECT 0.07 1.175 0.325 1.435 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3704 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.27 1.56 8.51 2.25 ;
        RECT 8.39 0.36 8.51 2.25 ;
        RECT 8.135 0.65 8.51 0.8 ;
        RECT 8.27 0.36 8.51 0.8 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.73 -0.18 7.97 0.32 ;
        RECT 7.79 -0.18 7.91 0.67 ;
        RECT 1.865 -0.18 2.105 0.32 ;
        RECT 0.685 -0.18 0.925 0.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.73 2.29 7.97 2.79 ;
        RECT 7.79 1.69 7.91 2.79 ;
        RECT 1.865 2.27 2.105 2.79 ;
        RECT 0.685 2.29 0.925 2.79 ;
        RECT 0.745 1.97 0.865 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.23 1.315 7.67 1.315 7.67 2.17 6.26 2.17 6.26 1.89 6.56 1.89 6.56 2.05 7.55 2.05 7.55 0.62 7.42 0.62 7.42 0.48 6.26 0.48 6.26 0.36 7.54 0.36 7.54 0.5 7.67 0.5 7.67 1.195 7.99 1.195 7.99 1.075 8.23 1.075 ;
      POLYGON 7.43 0.86 7.345 0.86 7.345 1.81 7.43 1.81 7.43 1.93 7.19 1.93 7.19 1.81 7.225 1.81 7.225 0.86 7.19 0.86 7.19 0.74 7.43 0.74 ;
      POLYGON 7.05 1.77 7.04 1.77 7.04 1.79 6.8 1.79 6.8 1.77 4.275 1.77 4.275 1.65 5.095 1.65 5.095 0.72 4.27 0.72 4.27 0.6 5.215 0.6 5.215 1.65 6.93 1.65 6.93 0.72 6.8 0.72 6.8 0.6 7.05 0.6 ;
      POLYGON 5.96 0.705 5.9 0.705 5.9 0.72 5.48 0.72 5.48 1.405 5.96 1.405 5.96 1.525 5.36 1.525 5.36 0.6 5.72 0.6 5.72 0.585 5.96 0.585 ;
      RECT 2.985 1.89 5.96 2.01 ;
      RECT 2.405 0.36 5.555 0.48 ;
      RECT 2.405 2.13 5.555 2.25 ;
      POLYGON 4.84 1.04 4.17 1.04 4.17 1.415 4.05 1.415 4.05 0.92 4.84 0.92 ;
      POLYGON 3.985 0.72 3.84 0.72 3.84 1.77 1.725 1.77 1.725 2.17 0.985 2.17 0.985 1.81 0.325 1.81 0.325 1.93 0.145 1.93 0.145 1.69 0.505 1.69 0.505 0.92 0.205 0.92 0.205 0.44 1.605 0.44 1.605 0.32 1.725 0.32 1.725 0.56 0.325 0.56 0.325 0.8 0.625 0.8 0.625 1.69 1.105 1.69 1.105 2.05 1.605 2.05 1.605 1.65 3.72 1.65 3.72 0.6 3.985 0.6 ;
      POLYGON 3.585 1.04 3.405 1.04 3.405 1 2.81 1 2.81 1.16 2.885 1.16 2.885 1.28 2.645 1.28 2.645 1.16 2.69 1.16 2.69 0.88 3.405 0.88 3.405 0.8 3.585 0.8 ;
      POLYGON 3.225 1.53 1.94 1.53 1.94 0.6 3.205 0.6 3.205 0.72 2.06 0.72 2.06 1.41 3.225 1.41 ;
      POLYGON 1.485 1.46 1.405 1.46 1.405 1.81 1.465 1.81 1.465 1.93 1.225 1.93 1.225 1.81 1.285 1.81 1.285 1.46 1.245 1.46 1.245 1.34 1.285 1.34 1.285 0.8 1.225 0.8 1.225 0.68 1.465 0.68 1.465 0.8 1.405 0.8 1.405 1.34 1.485 1.34 ;
  END
END XNOR3XL

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.09 0.29 1.42 ;
        RECT 0.07 1.105 0.22 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.08 0.835 1.47 ;
        RECT 0.65 1.08 0.835 1.46 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.355 0.885 1.67 1.145 ;
        RECT 1.355 0.67 1.475 2.07 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 1.775 -0.18 1.895 0.72 ;
        RECT 0.935 -0.18 1.055 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 1.42 1.895 2.79 ;
        RECT 0.935 1.59 1.055 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.195 1.23 1.075 1.23 1.075 0.96 0.53 0.96 0.53 1.59 0.635 1.59 0.635 1.83 0.515 1.83 0.515 1.71 0.41 1.71 0.41 0.96 0.235 0.96 0.235 0.67 0.355 0.67 0.355 0.84 1.195 0.84 ;
  END
END AND2X2

MACRO OR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 0.51 1.455 ;
        RECT 0.36 1 0.48 1.48 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1.02 0.815 1.455 ;
        RECT 0.65 1.02 0.815 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.205 1.435 1.42 ;
        RECT 1.175 1.04 1.295 1.42 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.655 1.295 1.96 1.435 ;
        RECT 1.81 1.175 1.96 1.435 ;
        RECT 1.815 0.4 1.935 0.64 ;
        RECT 1.81 0.52 1.93 1.435 ;
        RECT 1.655 1.295 1.775 1.66 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.235 1.54 1.355 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.615 1.04 1.495 1.04 1.495 0.92 1.055 0.92 1.055 1.72 0.155 1.72 0.155 1.6 0.935 1.6 0.935 0.88 0.135 0.88 0.135 0.4 0.255 0.4 0.255 0.76 0.975 0.76 0.975 0.4 1.095 0.4 1.095 0.8 1.615 0.8 ;
  END
END OR3XL

MACRO CLKBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX4 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.955 1.24 2.075 1.48 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.84 1.36 2.075 1.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.335 0.71 1.575 0.83 ;
        RECT 1.395 1.32 1.515 2.21 ;
        RECT 0.515 0.76 1.455 0.88 ;
        RECT 0.515 1.32 1.515 1.44 ;
        RECT 0.555 1.32 0.8 1.725 ;
        RECT 0.555 1.32 0.675 2.21 ;
        RECT 0.555 0.64 0.675 0.88 ;
        RECT 0.515 0.76 0.635 1.44 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.815 -0.18 1.935 0.7 ;
        RECT 0.915 0.52 1.155 0.64 ;
        RECT 0.915 -0.18 1.035 0.64 ;
        RECT 0.135 -0.18 0.255 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.815 1.845 1.935 2.79 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.355 2.21 2.235 2.21 2.235 1.12 1.415 1.12 1.415 1.17 1.175 1.17 1.175 1.12 0.995 1.12 0.995 1.17 0.755 1.17 0.755 1.05 0.875 1.05 0.875 1 2.235 1 2.235 0.65 2.355 0.65 ;
  END
END CLKBUFX4

MACRO AO22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X1 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.935 0.91 1.055 1.15 ;
        RECT 0.65 0.91 1.055 1.03 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.94 1.435 1.15 ;
        RECT 1.275 0.94 1.395 1.305 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.03 0.415 1.37 ;
        RECT 0.295 0.95 0.415 1.37 ;
        RECT 0.07 1.03 0.22 1.44 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 1.015 1.96 1.435 ;
        RECT 1.795 1 1.915 1.44 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.645 1.145 2.765 2.21 ;
        RECT 2.42 1.145 2.765 1.265 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.375 0.59 2.495 1.025 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.955 -0.18 2.075 0.64 ;
        RECT 0.41 -0.18 0.53 0.83 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.165 2.01 2.405 2.15 ;
        RECT 2.165 2.01 2.285 2.79 ;
        RECT 0.615 2.08 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.255 1.15 2.135 1.15 2.135 0.88 1.675 0.88 1.675 1.62 1.435 1.62 1.435 1.5 1.555 1.5 1.555 0.77 1.015 0.77 1.015 0.65 1.675 0.65 1.675 0.76 2.255 0.76 ;
      POLYGON 2.035 1.86 1.075 1.86 1.075 1.68 0.075 1.68 0.075 1.56 1.195 1.56 1.195 1.74 1.915 1.74 1.915 1.56 2.035 1.56 ;
  END
END AO22X1

MACRO NOR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.09 1.67 1.575 ;
        RECT 1.52 1.09 1.67 1.545 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.305 1.38 1.725 ;
        RECT 1.23 1.09 1.35 1.725 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 1.03 1.33 ;
        RECT 0.91 1.09 1.03 1.33 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.865 0.51 1.34 ;
        RECT 0.07 0.865 0.51 0.985 ;
        RECT 0.07 0.85 0.22 1.3 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4572 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 0.885 1.96 1.145 ;
        RECT 1.79 0.85 1.91 2.205 ;
        RECT 0.65 0.85 1.91 0.97 ;
        RECT 1.49 0.68 1.61 0.97 ;
        RECT 0.65 0.68 0.77 0.97 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.91 -0.18 2.03 0.73 ;
        RECT 1.07 -0.18 1.19 0.73 ;
        RECT 0.23 -0.18 0.35 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 0.43 1.555 0.55 2.79 ;
    END
  END VDD
END NOR4X1

MACRO DFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX4 0 0 ;
  SIZE 11.31 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 1.43 0.405 1.55 ;
        RECT 0.285 1.125 0.405 1.55 ;
        RECT 0.07 1.43 0.22 1.84 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.02 1.665 1.14 ;
        RECT 1.23 1.175 1.38 1.435 ;
        RECT 1.26 1.02 1.38 1.435 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 0.93 6.695 1.05 ;
        RECT 5.535 0.63 5.655 1.09 ;
        RECT 5.035 0.63 5.655 0.75 ;
        RECT 5.035 0.38 5.155 0.75 ;
        RECT 3.955 0.38 5.155 0.5 ;
        RECT 3.085 1.24 4.075 1.36 ;
        RECT 3.955 0.38 4.075 1.36 ;
        RECT 3.925 0.94 4.075 1.36 ;
        RECT 3.785 0.94 4.075 1.09 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.155 0.68 8.355 0.8 ;
        RECT 8.175 1.32 8.295 2.21 ;
        RECT 7.32 1.32 8.295 1.44 ;
        RECT 7.32 1.175 7.47 1.44 ;
        RECT 7.32 0.68 7.44 1.56 ;
        RECT 7.215 1.44 7.335 2.21 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.075 0.68 10.275 0.8 ;
        RECT 9.895 1.54 10.015 2.21 ;
        RECT 9.855 1.32 9.975 1.66 ;
        RECT 9.06 1.32 9.975 1.44 ;
        RECT 9.09 0.68 9.21 1.56 ;
        RECT 9.055 1.44 9.175 2.21 ;
        RECT 9.06 1.175 9.21 1.56 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.31 0.18 ;
        RECT 10.635 -0.18 10.755 0.67 ;
        RECT 9.555 -0.18 9.795 0.32 ;
        RECT 8.595 -0.18 8.835 0.32 ;
        RECT 7.635 -0.18 7.875 0.32 ;
        RECT 6.675 -0.18 6.915 0.32 ;
        RECT 5.275 0.39 5.515 0.51 ;
        RECT 5.395 -0.18 5.515 0.51 ;
        RECT 3.595 0.68 3.835 0.8 ;
        RECT 3.715 -0.18 3.835 0.8 ;
        RECT 1.685 0.54 1.925 0.66 ;
        RECT 1.685 -0.18 1.805 0.66 ;
        RECT 1.295 0.54 1.535 0.66 ;
        RECT 1.295 -0.18 1.415 0.66 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.31 2.79 ;
        RECT 10.315 1.56 10.435 2.79 ;
        RECT 9.475 1.56 9.595 2.79 ;
        RECT 8.635 1.56 8.755 2.79 ;
        RECT 7.755 1.56 7.875 2.79 ;
        RECT 6.795 1.73 6.915 2.79 ;
        RECT 5.955 1.73 6.075 2.79 ;
        RECT 5.115 1.73 5.235 2.79 ;
        RECT 3.735 2.29 3.975 2.79 ;
        RECT 2.535 2.2 2.775 2.79 ;
        RECT 1.285 2.23 1.405 2.79 ;
        RECT 0.135 1.97 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.175 0.86 10.995 0.86 10.995 1.42 10.855 1.42 10.855 2.21 10.735 2.21 10.735 1.42 10.095 1.42 10.095 1.28 10.335 1.28 10.335 1.3 10.875 1.3 10.875 0.74 11.055 0.74 11.055 0.62 11.175 0.62 ;
      POLYGON 10.715 1.18 10.595 1.18 10.595 0.91 10.395 0.91 10.395 0.56 8.595 0.56 8.595 1.08 8.555 1.08 8.555 1.2 8.435 1.2 8.435 0.96 8.475 0.96 8.475 0.56 6.215 0.56 6.215 0.61 5.975 0.61 5.975 0.49 6.095 0.49 6.095 0.44 10.515 0.44 10.515 0.79 10.715 0.79 ;
      POLYGON 7.055 1.61 6.495 1.61 6.495 2.21 6.375 2.21 6.375 1.61 5.655 1.61 5.655 2.21 5.535 2.21 5.535 1.61 5.055 1.61 5.055 1.55 4.935 1.55 4.935 1.43 5.175 1.43 5.175 1.49 6.935 1.49 6.935 1.24 7.055 1.24 ;
      POLYGON 5.915 1.37 5.295 1.37 5.295 0.99 4.575 0.99 4.575 1.97 4.455 1.97 4.455 0.75 4.615 0.75 4.615 0.62 4.735 0.62 4.735 0.87 5.415 0.87 5.415 1.25 5.915 1.25 ;
      POLYGON 4.935 1.23 4.815 1.23 4.815 2.21 4.375 2.21 4.375 2.23 4.135 2.23 4.135 2.21 4.095 2.21 4.095 2.17 3.615 2.17 3.615 2.25 2.895 2.25 2.895 2.08 2.39 2.08 2.39 2.22 2.15 2.22 2.15 2.11 1.065 2.11 1.065 2.25 0.945 2.25 0.945 2.11 0.675 2.11 0.675 2.2 0.555 2.2 0.555 2.08 0.545 2.08 0.545 0.68 0.665 0.68 0.665 1.96 0.675 1.96 0.675 1.99 2.005 1.99 2.005 1.96 3.015 1.96 3.015 2.13 3.495 2.13 3.495 2.05 4.215 2.05 4.215 2.09 4.695 2.09 4.695 1.11 4.935 1.11 ;
      POLYGON 4.315 1.72 4.155 1.72 4.155 1.85 4.035 1.85 4.035 1.6 2.765 1.6 2.765 1.48 4.195 1.48 4.195 0.62 4.315 0.62 ;
      POLYGON 3.665 1.12 2.505 1.12 2.505 1.48 2.285 1.48 2.285 1.7 2.105 1.7 2.105 1.84 1.985 1.84 1.985 1.58 2.165 1.58 2.165 1.36 2.385 1.36 2.385 0.68 2.625 0.68 2.625 0.8 2.505 0.8 2.505 1 3.665 1 ;
      POLYGON 3.595 0.48 2.165 0.48 2.165 0.9 1.905 0.9 1.905 1.34 2.025 1.34 2.025 1.46 1.785 1.46 1.785 0.9 1.055 0.9 1.055 1.69 0.985 1.69 0.985 1.81 0.865 1.81 0.865 1.57 0.935 1.57 0.935 0.48 1.055 0.48 1.055 0.78 2.045 0.78 2.045 0.36 3.595 0.36 ;
      POLYGON 3.375 2.01 3.135 2.01 3.135 1.84 2.405 1.84 2.405 1.6 2.525 1.6 2.525 1.72 3.255 1.72 3.255 1.89 3.375 1.89 ;
  END
END DFFRX4

MACRO AND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X4 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.72 0.51 1.2 ;
        RECT 0.36 0.72 0.51 1.175 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 0.96 0.99 1.2 ;
        RECT 0.65 0.96 0.99 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.35 1.36 1.64 1.48 ;
        RECT 1.35 1.24 1.47 1.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.79 0.885 3.12 1.145 ;
        RECT 1.91 1.32 2.91 1.44 ;
        RECT 2.79 0.67 2.91 1.44 ;
        RECT 2.75 1.32 2.87 2.21 ;
        RECT 1.83 0.72 2.91 0.84 ;
        RECT 2.55 0.67 2.91 0.84 ;
        RECT 1.91 1.32 2.03 2.21 ;
        RECT 1.71 0.67 1.95 0.79 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 3.03 -0.18 3.15 0.66 ;
        RECT 2.13 0.48 2.37 0.6 ;
        RECT 2.13 -0.18 2.25 0.6 ;
        RECT 1.35 -0.18 1.47 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 3.17 1.56 3.29 2.79 ;
        RECT 2.33 1.56 2.45 2.79 ;
        RECT 1.49 1.845 1.61 2.79 ;
        RECT 0.65 1.56 0.77 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.67 1.13 2.43 1.13 2.43 1.12 2.21 1.12 2.21 1.13 1.97 1.13 1.97 1.12 1.23 1.12 1.23 1.44 1.19 1.44 1.19 2.21 1.07 2.21 1.07 1.44 0.35 1.44 0.35 2.21 0.23 2.21 0.23 1.32 1.11 1.32 1.11 0.6 0.33 0.6 0.33 0.48 1.23 0.48 1.23 1 2.55 1 2.55 1.01 2.67 1.01 ;
  END
END AND3X4

MACRO SDFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX1 0 0 ;
  SIZE 13.05 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.905 1.21 2.145 1.385 ;
        RECT 1.755 1.23 2.015 1.43 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.735 2.13 7.575 2.25 ;
        RECT 6.735 1.8 6.855 2.25 ;
        RECT 5.105 1.8 6.855 1.92 ;
        RECT 5.105 1.4 5.225 1.92 ;
        RECT 3.635 1.4 5.225 1.52 ;
        RECT 3.635 1.23 3.755 1.52 ;
        RECT 3.335 1.27 3.755 1.39 ;
        RECT 3.495 1.23 3.755 1.39 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.56 1.03 10.68 1.465 ;
        RECT 10.51 1.03 10.68 1.445 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.8 1.465 11.025 1.77 ;
        RECT 10.83 1.455 11.025 1.77 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 1.4 12.455 1.67 ;
        RECT 12.19 1.4 12.455 1.65 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.95 1.16 12.75 1.28 ;
        RECT 12.195 0.94 12.455 1.28 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 1.295 1.485 2.14 ;
        RECT 1.365 0.61 1.485 0.85 ;
        RECT 1.23 1.175 1.425 1.435 ;
        RECT 1.305 0.73 1.425 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.05 0.18 ;
        RECT 12.19 -0.18 12.31 0.73 ;
        RECT 10.85 0.55 11.09 0.67 ;
        RECT 10.97 -0.18 11.09 0.67 ;
        RECT 9.65 -0.18 9.89 0.34 ;
        RECT 7.815 -0.18 7.935 0.86 ;
        RECT 3.015 -0.18 3.135 0.38 ;
        RECT 1.785 -0.18 1.905 0.85 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.05 2.79 ;
        RECT 12.305 2.03 12.545 2.15 ;
        RECT 12.305 2.03 12.425 2.79 ;
        RECT 10.865 1.95 10.985 2.79 ;
        RECT 9.885 1.6 10.005 2.79 ;
        RECT 7.695 2.13 7.935 2.25 ;
        RECT 7.695 2.13 7.815 2.79 ;
        RECT 6.035 2.29 6.275 2.79 ;
        RECT 4.355 2.12 4.595 2.24 ;
        RECT 4.355 2.12 4.475 2.79 ;
        RECT 3.075 1.75 3.195 2.79 ;
        RECT 1.785 1.55 1.905 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.99 1.97 12.905 1.97 12.905 2.09 12.785 2.09 12.785 1.91 11.925 1.91 11.925 2.25 11.145 2.25 11.145 1.03 11.59 1.03 11.59 1.15 11.265 1.15 11.265 2.13 11.805 2.13 11.805 1.51 11.925 1.51 11.925 1.79 12.87 1.79 12.87 0.73 12.73 0.73 12.73 0.49 12.85 0.49 12.85 0.61 12.99 0.61 ;
      POLYGON 11.83 1.39 11.685 1.39 11.685 2.01 11.445 2.01 11.445 1.27 11.71 1.27 11.71 0.73 11.405 0.73 11.405 0.91 10.61 0.91 10.61 0.48 10.13 0.48 10.13 0.58 9.6 0.58 9.6 0.62 8.995 0.62 8.995 0.74 9.275 0.74 9.275 1.89 9.195 1.89 9.195 2.01 9.075 2.01 9.075 1.77 9.155 1.77 9.155 0.86 8.875 0.86 8.875 0.5 9.48 0.5 9.48 0.46 10.01 0.46 10.01 0.36 10.73 0.36 10.73 0.79 11.285 0.79 11.285 0.61 11.55 0.61 11.55 0.49 11.67 0.49 11.67 0.61 11.83 0.61 ;
      POLYGON 10.49 0.72 10.39 0.72 10.39 1.565 10.44 1.565 10.44 2.07 10.32 2.07 10.32 1.685 10.27 1.685 10.27 1.22 9.835 1.22 9.835 1.34 9.715 1.34 9.715 1.1 10.27 1.1 10.27 0.72 10.25 0.72 10.25 0.6 10.49 0.6 ;
      POLYGON 9.635 0.86 9.585 0.86 9.585 2.25 8.835 2.25 8.835 2.22 8.235 2.22 8.235 2.01 6.975 2.01 6.975 1.68 6.755 1.68 6.755 1.56 6.365 1.56 6.365 1.23 6.485 1.23 6.485 1.44 6.875 1.44 6.875 1.56 7.095 1.56 7.095 1.89 8.235 1.89 8.235 1.48 8.435 1.48 8.435 1.72 8.355 1.72 8.355 2.1 8.835 2.1 8.835 1.12 8.795 1.12 8.795 1 9.035 1 9.035 1.12 8.955 1.12 8.955 2.13 9.465 2.13 9.465 0.86 9.395 0.86 9.395 0.74 9.635 0.74 ;
      POLYGON 8.715 1.98 8.475 1.98 8.475 1.86 8.555 1.86 8.555 1.2 7.235 1.2 7.235 0.96 7.355 0.96 7.355 1.08 8.555 1.08 8.555 0.86 8.455 0.86 8.455 0.62 8.575 0.62 8.575 0.74 8.675 0.74 8.675 1.86 8.715 1.86 ;
      POLYGON 8.115 1.44 7.335 1.44 7.335 1.65 7.455 1.65 7.455 1.77 7.215 1.77 7.215 1.44 6.995 1.44 6.995 1.11 6.245 1.11 6.245 1.64 5.765 1.64 5.765 1.52 6.125 1.52 6.125 1.02 5.865 1.02 5.865 0.62 5.985 0.62 5.985 0.9 6.245 0.9 6.245 0.99 6.975 0.99 6.975 0.62 7.095 0.62 7.095 0.99 7.115 0.99 7.115 1.32 8.115 1.32 ;
      POLYGON 7.575 0.8 7.335 0.8 7.335 0.5 6.855 0.5 6.855 0.68 6.735 0.68 6.735 0.8 6.495 0.8 6.495 0.68 6.615 0.68 6.615 0.56 6.735 0.56 6.735 0.38 7.455 0.38 7.455 0.68 7.575 0.68 ;
      POLYGON 6.615 2.17 4.715 2.17 4.715 2 4.23 2 4.23 2.13 4.235 2.13 4.235 2.25 3.995 2.25 3.995 2.12 3.315 2.12 3.315 1.63 2.955 1.63 2.955 2.11 2.265 2.11 2.265 1.91 2.205 1.91 2.205 1.67 2.265 1.67 2.265 0.61 2.385 0.61 2.385 1.99 2.835 1.99 2.835 1.51 3.435 1.51 3.435 2 4.11 2 4.11 1.88 4.835 1.88 4.835 2.05 6.615 2.05 ;
      POLYGON 6.005 1.38 5.885 1.38 5.885 1.26 5.625 1.26 5.625 0.48 5.185 0.48 5.185 0.36 5.745 0.36 5.745 1.14 6.005 1.14 ;
      POLYGON 5.585 1.64 5.345 1.64 5.345 1.52 5.385 1.52 5.385 1.28 3.915 1.28 3.915 1.11 3.035 1.11 3.035 1.24 2.915 1.24 2.915 0.99 4.035 0.99 4.035 1.16 5.385 1.16 5.385 0.62 5.505 0.62 5.505 1.52 5.585 1.52 ;
      POLYGON 5.085 0.92 4.995 0.92 4.995 1.04 4.155 1.04 4.155 0.62 4.275 0.62 4.275 0.92 4.875 0.92 4.875 0.8 4.965 0.8 4.965 0.62 5.085 0.62 ;
      POLYGON 4.985 1.76 3.675 1.76 3.675 1.88 3.555 1.88 3.555 1.64 4.985 1.64 ;
      POLYGON 4.755 0.8 4.515 0.8 4.515 0.5 4.035 0.5 4.035 0.72 3.735 0.72 3.735 0.8 3.495 0.8 3.495 0.68 3.615 0.68 3.615 0.6 3.915 0.6 3.915 0.38 4.635 0.38 4.635 0.68 4.755 0.68 ;
      POLYGON 3.795 0.48 3.375 0.48 3.375 0.75 3.11 0.75 3.11 0.87 2.775 0.87 2.775 0.9 2.715 0.9 2.715 1.87 2.595 1.87 2.595 0.75 2.655 0.75 2.655 0.49 2.145 0.49 2.145 1.09 1.785 1.09 1.785 1.11 1.545 1.11 1.545 0.97 2.025 0.97 2.025 0.37 2.775 0.37 2.775 0.75 2.99 0.75 2.99 0.63 3.255 0.63 3.255 0.36 3.795 0.36 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END SDFFNSRX1

MACRO DFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX1 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.565 0.96 6.945 1.21 ;
        RECT 6.685 0.94 6.945 1.21 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 1.155 0.995 1.32 ;
        RECT 0.595 1.185 0.855 1.38 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.215 1.22 2.595 1.4 ;
        RECT 2.335 1.195 2.595 1.4 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 1.34 0.255 1.99 ;
        RECT 0.135 0.555 0.255 0.795 ;
        RECT 0.07 1.175 0.235 1.435 ;
        RECT 0.115 0.675 0.235 1.46 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.035 0.46 7.275 0.58 ;
        RECT 7.035 -0.18 7.155 0.58 ;
        RECT 6.355 0.46 6.595 0.58 ;
        RECT 6.355 -0.18 6.475 0.58 ;
        RECT 4.495 -0.18 4.735 0.39 ;
        RECT 2.075 0.46 2.315 0.58 ;
        RECT 2.195 -0.18 2.315 0.58 ;
        RECT 0.495 0.675 0.735 0.795 ;
        RECT 0.495 -0.18 0.615 0.795 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.035 2.17 7.155 2.79 ;
        RECT 5.375 2.12 5.495 2.79 ;
        RECT 5.255 2.12 5.495 2.24 ;
        RECT 4.135 1.71 4.375 1.93 ;
        RECT 4.135 1.71 4.255 2.79 ;
        RECT 2.565 1.76 2.685 2.79 ;
        RECT 2.445 1.76 2.685 1.93 ;
        RECT 1.435 1.68 1.555 2.79 ;
        RECT 0.555 1.5 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.635 1.81 7.515 1.81 7.515 1.45 6.615 1.45 6.615 1.57 6.495 1.57 6.495 1.33 7.065 1.33 7.065 0.82 6.115 0.82 6.115 0.48 5.535 0.48 5.535 0.92 5.655 0.92 5.655 1.04 5.415 1.04 5.415 0.63 4.255 0.63 4.255 0.48 3.775 0.48 3.775 0.99 3.935 0.99 3.935 1.11 3.655 1.11 3.655 0.36 4.375 0.36 4.375 0.51 5.415 0.51 5.415 0.36 6.235 0.36 6.235 0.7 7.185 0.7 7.185 1.33 7.515 1.33 7.515 0.4 7.635 0.4 ;
      POLYGON 7.495 2.25 7.375 2.25 7.375 2.05 6.665 2.05 6.665 2.25 6.015 2.25 6.015 2 5.135 2 5.135 2.23 4.495 2.23 4.495 1.59 4.015 1.59 4.015 2.23 2.885 2.23 2.885 1.64 2.325 1.64 2.325 2.25 1.675 2.25 1.675 1.56 1.235 1.56 1.235 1.62 1.095 1.62 1.095 1.74 0.975 1.74 0.975 1.44 1.115 1.44 1.115 1.035 1.095 1.035 1.095 0.615 1.215 0.615 1.215 0.915 1.235 0.915 1.235 1.44 1.795 1.44 1.795 2.13 2.205 2.13 2.205 1.52 2.885 1.52 2.885 1.06 2.795 1.06 2.795 0.94 3.035 0.94 3.035 1.06 3.005 1.06 3.005 2.11 3.415 2.11 3.415 1.13 3.535 1.13 3.535 2.11 3.895 2.11 3.895 1.47 4.615 1.47 4.615 2.11 5.015 2.11 5.015 1.88 6.015 1.88 6.015 1.18 6.135 1.18 6.135 2.13 6.545 2.13 6.545 1.93 7.495 1.93 ;
      POLYGON 6.375 2.01 6.255 2.01 6.255 1.06 5.895 1.06 5.895 1.28 4.415 1.28 4.415 1.35 4.295 1.35 4.295 1.11 4.415 1.11 4.415 1.16 5.775 1.16 5.775 0.72 5.655 0.72 5.655 0.6 5.895 0.6 5.895 0.94 6.375 0.94 ;
      POLYGON 5.895 1.76 4.895 1.76 4.895 1.99 4.775 1.99 4.775 1.64 5.775 1.64 5.775 1.52 5.895 1.52 ;
      POLYGON 5.295 1.04 5.055 1.04 5.055 0.99 4.175 0.99 4.175 1.35 3.775 1.35 3.775 1.99 3.655 1.99 3.655 1.23 4.055 1.23 4.055 0.87 3.895 0.87 3.895 0.6 4.135 0.6 4.135 0.75 4.175 0.75 4.175 0.87 5.175 0.87 5.175 0.92 5.295 0.92 ;
      POLYGON 3.295 1.99 3.175 1.99 3.175 0.82 1.855 0.82 1.855 1.08 1.655 1.08 1.655 0.84 1.735 0.84 1.735 0.7 3.175 0.7 3.175 0.5 3.295 0.5 ;
      POLYGON 2.675 1.06 2.095 1.06 2.095 1.4 2.035 1.4 2.035 2.01 1.915 2.01 1.915 1.32 1.415 1.32 1.415 0.495 0.975 0.495 0.975 1.035 0.475 1.035 0.475 1.22 0.355 1.22 0.355 0.915 0.855 0.915 0.855 0.375 1.615 0.375 1.615 0.72 1.535 0.72 1.535 1.2 1.975 1.2 1.975 0.94 2.675 0.94 ;
  END
END DFFRHQX1

MACRO AOI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211XL 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.33 1.055 1.475 1.295 ;
        RECT 1.23 1.175 1.4 1.435 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 1.055 1.11 1.26 ;
        RECT 0.94 1.055 1.09 1.45 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.16 0.75 1.29 ;
        RECT 0.36 1.16 0.51 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.89 0.24 1.35 ;
        RECT 0.07 0.885 0.22 1.32 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.615 0.515 1.735 1.93 ;
        RECT 1.52 1.465 1.735 1.725 ;
        RECT 0.775 0.815 1.735 0.935 ;
        RECT 0.775 0.515 0.895 0.935 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 1.135 0.575 1.375 0.695 ;
        RECT 1.135 -0.18 1.255 0.695 ;
        RECT 0.135 -0.18 0.255 0.755 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 0.555 1.81 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.155 1.87 0.915 1.87 0.915 1.69 0.315 1.69 0.315 1.87 0.075 1.87 0.075 1.75 0.195 1.75 0.195 1.57 1.035 1.57 1.035 1.75 1.155 1.75 ;
  END
END AOI211XL

MACRO DFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX2 0 0 ;
  SIZE 8.7 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.45 0.855 1.68 ;
        RECT 0.715 1.16 0.835 1.68 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.475 1.27 2.715 1.44 ;
        RECT 2.335 1.23 2.595 1.43 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 1.45 6.075 1.67 ;
        RECT 5.825 1.28 5.945 1.67 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.715 1.465 6.89 1.725 ;
        RECT 6.715 0.8 6.835 2.15 ;
        RECT 6.525 0.8 6.835 0.92 ;
        RECT 6.525 0.68 6.645 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 1.465 7.76 1.725 ;
        RECT 7.555 1.465 7.675 2.15 ;
        RECT 7.425 0.74 7.665 0.86 ;
        RECT 7.465 0.74 7.585 1.62 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.7 0.18 ;
        RECT 7.905 -0.18 8.145 0.32 ;
        RECT 6.945 -0.18 7.185 0.32 ;
        RECT 6.045 -0.18 6.165 0.92 ;
        RECT 4.225 -0.18 4.345 0.86 ;
        RECT 2.505 0.51 2.745 0.63 ;
        RECT 2.505 -0.18 2.625 0.63 ;
        RECT 0.945 0.68 1.185 0.8 ;
        RECT 0.945 -0.18 1.065 0.8 ;
        RECT 0.555 -0.18 0.675 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.7 2.79 ;
        RECT 7.975 1.5 8.095 2.79 ;
        RECT 7.135 1.5 7.255 2.79 ;
        RECT 6.295 1.79 6.415 2.79 ;
        RECT 5.485 2.08 5.605 2.79 ;
        RECT 4.525 2.08 4.645 2.79 ;
        RECT 2.925 2.04 3.045 2.79 ;
        RECT 1.845 2.29 2.085 2.79 ;
        RECT 0.615 2.12 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.565 1.345 8.515 1.345 8.515 1.74 8.395 1.74 8.395 1.345 7.705 1.345 7.705 1.225 8.445 1.225 8.445 0.68 8.565 0.68 ;
      POLYGON 8.505 0.52 8.385 0.52 8.385 0.56 7.075 0.56 7.075 1.26 6.955 1.26 6.955 0.56 6.405 0.56 6.405 1.24 6.285 1.24 6.285 1.16 5.805 1.16 5.805 0.56 5.285 0.56 5.285 0.68 5.445 0.68 5.445 1.36 5.125 1.36 5.125 1.72 5.005 1.72 5.005 1.36 4.505 1.36 4.505 1.34 4.385 1.34 4.385 1.22 4.625 1.22 4.625 1.24 5.325 1.24 5.325 0.8 5.165 0.8 5.165 0.44 5.925 0.44 5.925 1.04 6.285 1.04 6.285 0.44 8.265 0.44 8.265 0.4 8.505 0.4 ;
      POLYGON 5.995 2.03 5.875 2.03 5.875 1.96 4.405 1.96 4.405 2.23 3.865 2.23 3.865 2.25 3.625 2.25 3.625 2.23 3.165 2.23 3.165 1.92 2.805 1.92 2.805 2.17 1.385 2.17 1.385 2.1 0.855 2.1 0.855 2 0.395 2 0.395 2.16 0.275 2.16 0.275 1.88 0.975 1.88 0.975 1.98 1.625 1.98 1.625 2.05 2.685 2.05 2.685 1.8 3.285 1.8 3.285 2.11 4.285 2.11 4.285 1.84 5.565 1.84 5.565 0.68 5.685 0.68 5.685 1.79 5.995 1.79 ;
      POLYGON 5.205 1.12 4.965 1.12 4.965 1.1 4.265 1.1 4.265 1.72 4.005 1.72 4.005 1.81 3.765 1.81 3.765 1.69 3.885 1.69 3.885 1.6 4.145 1.6 4.145 1.1 3.585 1.1 3.585 0.62 3.705 0.62 3.705 0.98 5.085 0.98 5.085 1 5.205 1 ;
      POLYGON 4.025 1.48 3.905 1.48 3.905 1.36 3.345 1.36 3.345 0.5 2.985 0.5 2.985 0.87 2.265 0.87 2.265 0.56 1.425 0.56 1.425 1.04 1.195 1.04 1.195 1.4 1.075 1.4 1.075 1.04 0.255 1.04 0.255 1.72 0.135 1.72 0.135 0.74 0.075 0.74 0.075 0.62 0.315 0.62 0.315 0.74 0.255 0.74 0.255 0.92 1.305 0.92 1.305 0.44 1.725 0.44 1.725 0.36 1.965 0.36 1.965 0.44 2.385 0.44 2.385 0.75 2.865 0.75 2.865 0.38 3.465 0.38 3.465 1.24 4.025 1.24 ;
      POLYGON 3.525 1.99 3.405 1.99 3.405 1.68 2.095 1.68 2.095 1.41 2.215 1.41 2.215 1.56 3.105 1.56 3.105 0.62 3.225 0.62 3.225 1.56 3.525 1.56 ;
      POLYGON 2.985 1.12 2.715 1.12 2.715 1.11 1.705 1.11 1.705 1.48 1.515 1.48 1.515 1.64 1.335 1.64 1.335 1.76 1.215 1.76 1.215 1.52 1.395 1.52 1.395 1.36 1.585 1.36 1.585 0.68 1.825 0.68 1.825 0.8 1.705 0.8 1.705 0.99 2.835 0.99 2.835 1 2.985 1 ;
      POLYGON 2.565 1.93 2.06 1.93 2.06 1.92 1.795 1.92 1.795 1.86 1.635 1.86 1.635 1.6 1.755 1.6 1.755 1.74 1.915 1.74 1.915 1.8 2.18 1.8 2.18 1.81 2.565 1.81 ;
  END
END DFFRX2

MACRO AND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X6 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.84 0.97 2.08 1.09 ;
        RECT 1.84 0.595 1.96 1.09 ;
        RECT 1.81 0.595 1.96 0.855 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.09 ;
        RECT 1.3 1.21 2.78 1.33 ;
        RECT 2.66 0.94 2.78 1.33 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.45 3.3 1.57 ;
        RECT 3.18 1.22 3.3 1.57 ;
        RECT 0.94 1.175 1.09 1.57 ;
        RECT 0.76 1.28 1.09 1.4 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.5 1.465 3.7 1.725 ;
        RECT 0.5 1.69 3.67 1.81 ;
        RECT 3.5 1.22 3.62 1.81 ;
        RECT 0.5 1.22 0.62 1.81 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.08 1.41 6.2 2.21 ;
        RECT 4.4 1.41 6.2 1.53 ;
        RECT 5.64 0.795 5.94 0.915 ;
        RECT 5.82 0.4 5.94 0.915 ;
        RECT 4.08 0.93 5.76 1.05 ;
        RECT 5.64 0.795 5.76 1.05 ;
        RECT 5.24 1.41 5.36 2.21 ;
        RECT 5 1.175 5.15 1.53 ;
        RECT 5 0.93 5.12 1.53 ;
        RECT 4.98 0.4 5.1 1.05 ;
        RECT 4.4 1.41 4.52 2.21 ;
        RECT 4.08 0.4 4.2 1.05 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.4 -0.18 5.52 0.81 ;
        RECT 4.56 -0.18 4.68 0.81 ;
        RECT 3.6 0.46 3.84 0.58 ;
        RECT 3.6 -0.18 3.72 0.58 ;
        RECT 0.34 -0.18 0.46 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.66 1.65 5.78 2.79 ;
        RECT 4.82 1.65 4.94 2.79 ;
        RECT 3.86 2.17 4.1 2.29 ;
        RECT 3.86 2.17 3.98 2.79 ;
        RECT 2.9 2.17 3.14 2.29 ;
        RECT 2.9 2.17 3.02 2.79 ;
        RECT 1.94 2.17 2.18 2.29 ;
        RECT 1.94 2.17 2.06 2.79 ;
        RECT 0.98 2.17 1.22 2.29 ;
        RECT 0.98 2.17 1.1 2.79 ;
        RECT 0.14 1.56 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.88 1.29 3.94 1.29 3.94 2.05 3.56 2.05 3.56 2.21 3.44 2.21 3.44 2.05 2.6 2.05 2.6 2.21 2.48 2.21 2.48 2.05 1.64 2.05 1.64 2.21 1.52 2.21 1.52 2.05 0.68 2.05 0.68 2.21 0.56 2.21 0.56 1.93 3.82 1.93 3.82 0.82 2.24 0.82 2.24 0.77 2.12 0.77 2.12 0.65 2.36 0.65 2.36 0.7 3.94 0.7 3.94 1.17 4.88 1.17 ;
  END
END AND4X6

MACRO OR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X4 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.95 0.51 1.19 ;
        RECT 0.07 0.95 0.51 1.07 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.45 1.09 1.725 ;
        RECT 0.93 1.355 1.06 1.475 ;
        RECT 0.93 1.22 1.05 1.475 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.39 0.74 2.51 1.68 ;
        RECT 2.35 1.56 2.47 2.21 ;
        RECT 1.51 1.32 2.51 1.44 ;
        RECT 1.57 0.74 2.51 0.86 ;
        RECT 2.35 0.62 2.47 0.86 ;
        RECT 1.45 0.69 1.69 0.81 ;
        RECT 1.51 1.32 1.63 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.77 -0.18 2.89 0.68 ;
        RECT 1.87 0.5 2.11 0.62 ;
        RECT 1.87 -0.18 1.99 0.62 ;
        RECT 1.09 -0.18 1.21 0.68 ;
        RECT 0.25 -0.18 0.37 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.77 1.56 2.89 2.79 ;
        RECT 1.93 1.56 2.05 2.79 ;
        RECT 1.09 1.845 1.21 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.27 1.15 2.03 1.15 2.03 1.1 1.85 1.1 1.85 1.15 1.61 1.15 1.61 1.1 0.79 1.1 0.79 1.43 0.57 1.43 0.57 2.21 0.45 2.21 0.45 1.31 0.67 1.31 0.67 0.63 0.79 0.63 0.79 0.98 2.15 0.98 2.15 1.03 2.27 1.03 ;
  END
END OR2X4

MACRO NAND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 0.595 1.67 1.18 ;
        RECT 1.52 0.595 1.67 1.02 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.595 1.38 1 ;
        RECT 1.21 0.78 1.33 1.2 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.89 0.96 1.01 1.2 ;
        RECT 0.65 0.96 1.01 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 0.885 0.53 1.145 ;
        RECT 0.235 0.94 0.47 1.18 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5364 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 1.175 1.96 1.435 ;
        RECT 0.63 1.32 1.91 1.44 ;
        RECT 1.79 0.62 1.91 1.44 ;
        RECT 1.47 1.32 1.59 2.21 ;
        RECT 0.63 1.32 0.75 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 0.41 -0.18 0.53 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.89 1.56 2.01 2.79 ;
        RECT 1.05 1.56 1.17 2.79 ;
        RECT 0.21 1.56 0.33 2.79 ;
    END
  END VDD
END NAND4X1

MACRO NAND3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX4 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.575 0.97 3.815 1.09 ;
        RECT 3.575 0.82 3.695 1.09 ;
        RECT 2.2 0.82 3.695 0.94 ;
        RECT 1.615 0.97 2.32 1.09 ;
        RECT 2.2 0.82 2.32 1.09 ;
        RECT 1.755 0.94 2.015 1.09 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.085 0.985 5.415 1.12 ;
        RECT 4.945 0.94 5.205 1.105 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.935 1.08 4.675 1.2 ;
        RECT 3.235 1.21 4.055 1.33 ;
        RECT 3.935 1.08 4.055 1.33 ;
        RECT 3.235 1.06 3.355 1.33 ;
        RECT 2.44 1.06 3.355 1.18 ;
        RECT 1.115 1.21 2.56 1.33 ;
        RECT 2.44 1.06 2.56 1.33 ;
        RECT 1.115 1.08 1.235 1.33 ;
        RECT 0.885 0.94 1.145 1.2 ;
        RECT 0.755 1.08 1.235 1.2 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5232 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.755 1.56 4.875 2.21 ;
        RECT 0.255 1.69 4.875 1.81 ;
        RECT 3.915 1.69 4.035 2.21 ;
        RECT 0.255 0.58 3.895 0.7 ;
        RECT 3.075 1.69 3.195 2.21 ;
        RECT 2.235 1.69 2.355 2.21 ;
        RECT 1.395 1.69 1.515 2.21 ;
        RECT 0.555 1.56 0.675 2.21 ;
        RECT 0.07 1.465 0.375 1.725 ;
        RECT 0.255 0.58 0.375 1.81 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 4.975 -0.18 5.095 0.64 ;
        RECT 2.495 0.34 2.735 0.46 ;
        RECT 2.495 -0.18 2.615 0.46 ;
        RECT 0.215 0.34 0.455 0.46 ;
        RECT 0.215 -0.18 0.335 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.175 1.56 5.295 2.79 ;
        RECT 4.335 1.93 4.455 2.79 ;
        RECT 3.495 1.93 3.615 2.79 ;
        RECT 2.655 1.93 2.775 2.79 ;
        RECT 1.815 1.93 1.935 2.79 ;
        RECT 0.975 1.93 1.095 2.79 ;
        RECT 0.135 1.93 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.715 2.21 5.595 2.21 5.595 1.52 5.535 1.52 5.535 1.4 4.915 1.4 4.915 1.44 4.385 1.44 4.385 1.57 0.82 1.57 0.82 1.44 0.495 1.44 0.495 1.2 0.615 1.2 0.615 1.32 0.94 1.32 0.94 1.45 2.835 1.45 2.835 1.3 3.075 1.3 3.075 1.45 4.265 1.45 4.265 1.32 4.795 1.32 4.795 1.28 5.535 1.28 5.535 0.865 5.395 0.865 5.395 0.59 5.515 0.59 5.515 0.745 5.655 0.745 5.655 1.4 5.715 1.4 ;
  END
END NAND3BX4

MACRO SDFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX4 0 0 ;
  SIZE 16.24 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.675 0.36 1.795 1.41 ;
        RECT 1.015 0.36 1.795 0.48 ;
        RECT 1.015 0.96 1.235 1.2 ;
        RECT 0.375 0.935 1.135 1.055 ;
        RECT 1.015 0.36 1.135 1.2 ;
        RECT 0.94 0.595 1.135 1.055 ;
        RECT 0.375 0.935 0.495 1.175 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.895 1.485 ;
        RECT 0.65 1.175 0.8 1.49 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.145 2.25 1.435 ;
        RECT 1.995 0.99 2.115 1.265 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.095 2.54 1.47 ;
        RECT 2.39 0.96 2.51 1.47 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.155 0.97 6.275 1.21 ;
        RECT 5.815 0.97 6.275 1.09 ;
        RECT 5.815 0.94 6.075 1.09 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.535 1.09 7.415 1.21 ;
        RECT 6.395 0.94 6.655 1.09 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.835 0.74 13.035 0.86 ;
        RECT 12.735 1.42 12.855 2.19 ;
        RECT 12.555 1.42 12.855 1.54 ;
        RECT 11.96 1.3 12.675 1.42 ;
        RECT 11.96 1.175 12.11 1.435 ;
        RECT 11.96 0.74 12.08 1.54 ;
        RECT 11.895 1.42 12.015 2.19 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.755 0.74 14.955 0.86 ;
        RECT 14.415 1.42 14.535 2.19 ;
        RECT 14.235 1.42 14.535 1.54 ;
        RECT 13.7 1.3 14.355 1.42 ;
        RECT 13.575 1.42 13.875 1.54 ;
        RECT 13.755 0.74 13.875 1.54 ;
        RECT 13.7 1.175 13.875 1.54 ;
        RECT 13.575 1.42 13.695 2.19 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 16.24 0.18 ;
        RECT 15.315 -0.18 15.435 0.73 ;
        RECT 14.235 -0.18 14.475 0.38 ;
        RECT 13.275 -0.18 13.515 0.38 ;
        RECT 12.315 -0.18 12.555 0.38 ;
        RECT 11.355 -0.18 11.475 0.82 ;
        RECT 10.515 -0.18 10.635 0.86 ;
        RECT 7.015 0.61 7.255 0.73 ;
        RECT 7.135 -0.18 7.255 0.73 ;
        RECT 4.22 -0.18 4.46 0.32 ;
        RECT 1.915 -0.18 2.035 0.84 ;
        RECT 0.555 -0.18 0.675 0.815 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 16.24 2.79 ;
        RECT 14.835 1.54 14.955 2.79 ;
        RECT 13.995 1.54 14.115 2.79 ;
        RECT 13.155 1.54 13.275 2.79 ;
        RECT 12.315 1.54 12.435 2.79 ;
        RECT 11.475 1.64 11.595 2.79 ;
        RECT 10.635 1.7 10.755 2.79 ;
        RECT 9.515 1.88 9.755 2 ;
        RECT 9.515 1.88 9.635 2.79 ;
        RECT 6.375 2.13 6.615 2.25 ;
        RECT 6.375 2.13 6.495 2.79 ;
        RECT 4.835 2.2 5.075 2.79 ;
        RECT 4.22 2.17 4.34 2.79 ;
        RECT 4.1 2.17 4.34 2.29 ;
        RECT 2.145 2.23 2.265 2.79 ;
        RECT 0.675 1.85 0.795 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 15.855 0.92 15.695 0.92 15.695 1.42 15.375 1.42 15.375 2.19 15.255 2.19 15.255 1.42 14.655 1.42 14.655 1.28 14.895 1.28 14.895 1.3 15.575 1.3 15.575 0.8 15.735 0.8 15.735 0.68 15.855 0.68 ;
      POLYGON 15.455 1.18 15.215 1.18 15.215 0.97 15.075 0.97 15.075 0.62 11.715 0.62 11.715 1.06 11.215 1.06 11.215 1.28 11.775 1.28 11.775 1.4 11.215 1.4 11.215 1.76 11.175 1.76 11.175 2.16 11.055 2.16 11.055 1.64 11.095 1.64 11.095 1.24 9.975 1.24 9.975 1.12 10.935 1.12 10.935 0.68 11.055 0.68 11.055 0.94 11.595 0.94 11.595 0.5 15.195 0.5 15.195 0.85 15.335 0.85 15.335 1.06 15.455 1.06 ;
      POLYGON 10.975 1.52 8.505 1.52 8.505 1.77 8.385 1.77 8.385 0.87 8.365 0.87 8.365 0.63 8.485 0.63 8.485 0.75 8.505 0.75 8.505 1.4 10.735 1.4 10.735 1.36 10.975 1.36 ;
      POLYGON 10.395 1.88 9.875 1.88 9.875 1.76 8.745 1.76 8.745 1.64 9.995 1.64 9.995 1.76 10.395 1.76 ;
      POLYGON 10.215 0.86 10.095 0.86 10.095 0.56 9.435 0.56 9.435 0.8 9.195 0.8 9.195 0.68 9.315 0.68 9.315 0.44 10.215 0.44 ;
      POLYGON 9.855 0.8 9.675 0.8 9.675 1.04 8.865 1.04 8.865 0.63 8.985 0.63 8.985 0.92 9.555 0.92 9.555 0.68 9.855 0.68 ;
      POLYGON 9.595 1.28 8.625 1.28 8.625 0.51 7.685 0.51 7.685 0.74 7.675 0.74 7.675 1.41 7.695 1.41 7.695 1.53 7.455 1.53 7.455 1.41 7.555 1.41 7.555 0.97 6.775 0.97 6.775 0.48 6.195 0.48 6.195 0.36 6.895 0.36 6.895 0.85 7.375 0.85 7.375 0.62 7.565 0.62 7.565 0.39 8.745 0.39 8.745 1.16 9.595 1.16 ;
      POLYGON 9.325 2.05 9.085 2.05 9.085 2.01 6.975 2.01 6.975 1.77 5.675 1.77 5.675 1.57 4.98 1.57 4.98 1.33 5.1 1.33 5.1 1.45 5.795 1.45 5.795 1.65 7.095 1.65 7.095 1.89 8.145 1.89 8.145 1.23 8.085 1.23 8.085 0.99 8.205 0.99 8.205 1.11 8.265 1.11 8.265 1.89 9.205 1.89 9.205 1.93 9.325 1.93 ;
      POLYGON 8.305 2.25 6.735 2.25 6.735 2.01 5.435 2.01 5.435 1.81 4.58 1.81 4.58 1.69 4.7 1.69 4.7 1.44 3.74 1.44 3.74 1.56 3.62 1.56 3.62 1.32 4.715 1.32 4.715 0.84 4.635 0.84 4.635 0.72 4.875 0.72 4.875 0.84 4.835 0.84 4.835 1.44 4.82 1.44 4.82 1.69 5.555 1.69 5.555 1.89 6.855 1.89 6.855 2.13 8.305 2.13 ;
      POLYGON 8.065 0.87 7.965 0.87 7.965 1.53 8.025 1.53 8.025 1.77 7.215 1.77 7.215 1.53 5.915 1.53 5.915 1.33 5.575 1.33 5.575 1.1 4.995 1.1 4.995 0.56 3.98 0.56 3.98 0.48 3.86 0.48 3.86 0.36 4.1 0.36 4.1 0.44 5.115 0.44 5.115 0.98 5.575 0.98 5.575 0.68 5.835 0.68 5.835 0.8 5.695 0.8 5.695 1.21 6.035 1.21 6.035 1.41 7.335 1.41 7.335 1.65 7.845 1.65 7.845 0.75 7.945 0.75 7.945 0.63 8.065 0.63 ;
      POLYGON 6.255 0.8 5.955 0.8 5.955 0.56 5.455 0.56 5.455 0.62 5.355 0.62 5.355 0.86 5.235 0.86 5.235 0.5 5.335 0.5 5.335 0.44 6.075 0.44 6.075 0.68 6.255 0.68 ;
      POLYGON 5.92 2.25 5.195 2.25 5.195 2.05 3.4 2.05 3.4 1.8 3.38 1.8 3.38 0.62 3.5 0.62 3.5 1.68 3.52 1.68 3.52 1.93 5.315 1.93 5.315 2.13 5.92 2.13 ;
      POLYGON 4.595 1.16 3.8 1.16 3.8 1.2 3.68 1.2 3.68 1.16 3.62 1.16 3.62 0.5 3.26 0.5 3.26 1.56 3.14 1.56 3.14 0.5 2.595 0.5 2.595 0.72 2.78 0.72 2.78 1.71 2.71 1.71 2.71 1.83 2.59 1.83 2.59 1.59 2.66 1.59 2.66 0.84 2.475 0.84 2.475 0.38 3.74 0.38 3.74 0.96 3.8 0.96 3.8 1.04 4.595 1.04 ;
      POLYGON 3.1 2.07 1.415 2.07 1.415 0.84 1.255 0.84 1.255 0.6 1.375 0.6 1.375 0.72 1.535 0.72 1.535 1.95 2.98 1.95 2.98 1.83 2.9 1.83 2.9 0.62 3.02 0.62 3.02 1.71 3.1 1.71 ;
      POLYGON 1.295 1.73 0.375 1.73 0.375 1.97 0.255 1.97 0.255 1.85 0.135 1.85 0.135 0.575 0.255 0.575 0.255 1.61 1.175 1.61 1.175 1.41 1.295 1.41 ;
  END
END SDFFNSRX4

MACRO NAND2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BXL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.49 0.865 0.635 1.105 ;
        RECT 0.36 0.885 0.535 1.145 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.275 1.365 ;
        RECT 1.155 1.125 1.275 1.365 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.315 0.675 1.685 ;
        RECT 0.07 1.315 0.675 1.435 ;
        RECT 0.12 0.645 0.37 0.765 ;
        RECT 0.25 0.525 0.37 0.765 ;
        RECT 0.07 1.175 0.24 1.435 ;
        RECT 0.12 0.645 0.24 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.97 -0.18 1.09 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.005 2.085 1.125 2.79 ;
        RECT 0.135 1.565 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.605 1.685 1.485 1.685 1.485 1.565 1.395 1.565 1.395 1.005 1.035 1.005 1.035 1.045 0.755 1.045 0.755 0.925 0.915 0.925 0.915 0.885 1.395 0.885 1.395 0.765 1.39 0.765 1.39 0.525 1.51 0.525 1.51 0.645 1.515 0.645 1.515 1.445 1.605 1.445 ;
  END
END NAND2BXL

MACRO DFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX4 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 1 0.53 1.485 ;
        RECT 0.36 1 0.53 1.455 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 1 0.87 1.38 ;
        RECT 0.65 1.13 0.8 1.5 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.45 1.255 5.57 1.495 ;
        RECT 4.71 1.255 5.57 1.375 ;
        RECT 4.77 0.395 4.89 1.375 ;
        RECT 4.71 1.175 4.86 1.435 ;
        RECT 3.385 0.395 4.89 0.515 ;
        RECT 2.905 0.98 3.505 1.1 ;
        RECT 3.385 0.395 3.505 1.1 ;
        RECT 2.905 0.36 3.025 1.1 ;
        RECT 2.785 0.36 3.025 0.48 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.97 1.44 8.09 2.21 ;
        RECT 6.89 0.8 7.97 0.92 ;
        RECT 7.85 0.68 7.97 0.92 ;
        RECT 7.79 1.44 8.09 1.56 ;
        RECT 7.31 1.32 7.91 1.44 ;
        RECT 7.31 1.175 7.47 1.44 ;
        RECT 7.13 1.44 7.43 1.56 ;
        RECT 7.31 0.8 7.43 1.56 ;
        RECT 7.13 1.44 7.25 2.21 ;
        RECT 6.89 0.68 7.01 0.92 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.81 0.8 9.89 0.92 ;
        RECT 9.77 0.68 9.89 0.92 ;
        RECT 9.65 1.44 9.77 2.21 ;
        RECT 9.47 1.44 9.77 1.56 ;
        RECT 8.8 1.32 9.59 1.44 ;
        RECT 8.81 0.68 8.93 2.21 ;
        RECT 8.77 1.175 8.93 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.25 -0.18 10.37 0.73 ;
        RECT 9.23 -0.18 9.47 0.32 ;
        RECT 8.27 -0.18 8.51 0.32 ;
        RECT 7.31 -0.18 7.55 0.32 ;
        RECT 6.41 -0.18 6.53 0.82 ;
        RECT 5.57 -0.18 5.69 0.875 ;
        RECT 3.145 -0.18 3.265 0.86 ;
        RECT 1.995 -0.18 2.235 0.32 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.07 1.6 10.19 2.79 ;
        RECT 9.23 1.56 9.35 2.79 ;
        RECT 8.39 1.56 8.51 2.79 ;
        RECT 7.55 1.56 7.67 2.79 ;
        RECT 6.71 1.56 6.83 2.79 ;
        RECT 5.75 1.94 5.99 2.15 ;
        RECT 5.75 1.94 5.87 2.79 ;
        RECT 4.85 2.18 5.09 2.3 ;
        RECT 4.85 2.18 4.97 2.79 ;
        RECT 2.83 2.28 3.07 2.79 ;
        RECT 1.93 2.1 2.05 2.79 ;
        RECT 0.59 1.62 0.71 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.79 1.48 10.61 1.48 10.61 2.21 10.49 2.21 10.49 1.48 9.915 1.48 9.915 1.24 10.035 1.24 10.035 1.36 10.67 1.36 10.67 0.68 10.79 0.68 ;
      POLYGON 10.395 1.24 10.275 1.24 10.275 0.97 10.01 0.97 10.01 0.56 6.77 0.56 6.77 1.04 6.97 1.04 6.97 1.28 6.85 1.28 6.85 1.16 6.35 1.16 6.35 2.21 6.23 2.21 6.23 1.135 5.01 1.135 5.01 1.015 5.99 1.015 5.99 0.68 6.11 0.68 6.11 0.94 6.65 0.94 6.65 0.44 10.13 0.44 10.13 0.85 10.395 0.85 ;
      POLYGON 6.09 1.59 5.81 1.59 5.81 1.82 4.22 1.82 4.22 2.09 4.1 2.09 4.1 1.7 4.47 1.7 4.47 0.935 4.53 0.935 4.53 0.635 4.65 0.635 4.65 1.055 4.59 1.055 4.59 1.7 5.69 1.7 5.69 1.47 5.97 1.47 5.97 1.35 6.09 1.35 ;
      RECT 4.46 1.94 5.57 2.06 ;
      POLYGON 4.35 1.58 3.8 1.58 3.8 2.13 3.68 2.13 3.68 1.92 3.07 1.92 3.07 1.74 2.41 1.74 2.41 1.5 2.425 1.5 2.425 1.02 1.775 1.02 1.775 0.9 2.305 0.9 2.305 0.68 2.425 0.68 2.425 0.84 2.545 0.84 2.545 1.62 3.19 1.62 3.19 1.8 3.68 1.8 3.68 1.46 4.23 1.46 4.23 0.815 4.05 0.815 4.05 0.695 4.35 0.695 ;
      POLYGON 4.11 1.34 3.55 1.34 3.55 1.68 3.31 1.68 3.31 1.56 3.43 1.56 3.43 1.34 2.665 1.34 2.665 0.72 2.545 0.72 2.545 0.56 1.635 0.56 1.635 0.98 1.515 0.98 1.515 0.44 2.665 0.44 2.665 0.6 2.785 0.6 2.785 1.22 3.625 1.22 3.625 0.68 3.745 0.68 3.745 1.22 3.99 1.22 3.99 0.96 4.11 0.96 ;
      POLYGON 3.39 2.16 2.83 2.16 2.83 1.98 1.51 1.98 1.51 2.2 1.39 2.2 1.39 1.98 0.99 1.98 0.99 0.88 0.24 0.88 0.24 1.575 0.29 1.575 0.29 1.815 0.17 1.815 0.17 1.695 0.12 1.695 0.12 0.64 0.135 0.64 0.135 0.4 0.255 0.4 0.255 0.76 1.035 0.76 1.035 0.74 1.155 0.74 1.155 0.98 1.11 0.98 1.11 1.86 2.95 1.86 2.95 2.04 3.39 2.04 ;
      POLYGON 2.305 1.36 1.395 1.36 1.395 1.62 1.35 1.62 1.35 1.74 1.23 1.74 1.23 1.5 1.275 1.5 1.275 0.4 1.395 0.4 1.395 1.24 2.305 1.24 ;
  END
END DFFSX4

MACRO AND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X2 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.985 0.24 1.435 ;
        RECT 0.12 0.96 0.24 1.435 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.675 0.96 0.795 1.395 ;
        RECT 0.36 1.02 0.795 1.14 ;
        RECT 0.36 1.02 0.51 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.155 1.23 1.435 1.46 ;
        RECT 1.155 1.23 1.275 1.64 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.885 1.96 1.145 ;
        RECT 1.815 0.885 1.935 2.035 ;
        RECT 1.635 0.885 1.96 1.025 ;
        RECT 1.635 0.61 1.755 1.025 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 2.055 -0.18 2.175 0.66 ;
        RECT 1.215 -0.18 1.335 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 2.235 1.385 2.355 2.79 ;
        RECT 1.395 1.675 1.515 2.79 ;
        RECT 0.555 1.795 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.11 1.035 1.11 1.035 1.76 1.095 1.76 1.095 2 0.975 2 0.975 1.88 0.915 1.88 0.915 1.675 0.315 1.675 0.315 1.855 0.075 1.855 0.075 1.735 0.195 1.735 0.195 1.555 0.915 1.555 0.915 0.84 0.195 0.84 0.195 0.6 0.315 0.6 0.315 0.72 1.035 0.72 1.035 0.99 1.515 0.99 ;
  END
END AND3X2

MACRO ADDHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHXL 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.305 0.4 2.545 0.52 ;
        RECT 1.825 1.02 2.425 1.14 ;
        RECT 2.305 0.4 2.425 1.14 ;
        RECT 1.825 0.405 1.945 1.14 ;
        RECT 0.855 0.405 1.945 0.525 ;
        RECT 0.65 0.885 0.975 1.045 ;
        RECT 0.855 0.405 0.975 1.045 ;
        RECT 0.7 0.885 0.82 1.165 ;
        RECT 0.65 0.885 0.82 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.17 1.225 1.4 ;
        RECT 1.105 1.155 1.225 1.4 ;
        RECT 0.94 1.17 1.09 1.435 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.585 0.255 1.83 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.405 0.78 4.525 1.7 ;
        RECT 4.385 1.465 4.505 1.82 ;
        RECT 4.385 0.66 4.505 0.9 ;
        RECT 4.13 1.465 4.505 1.725 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 3.945 -0.18 4.065 0.38 ;
        RECT 2.065 -0.18 2.185 0.9 ;
        RECT 0.495 0.645 0.735 0.765 ;
        RECT 0.615 -0.18 0.735 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 3.945 2.22 4.065 2.79 ;
        RECT 2.105 1.76 2.345 1.88 ;
        RECT 2.105 1.76 2.225 2.79 ;
        RECT 1.455 2.09 1.575 2.79 ;
        RECT 0.615 2.23 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.285 1.18 3.825 1.18 3.825 1.66 3.425 1.66 3.425 1.76 3.185 1.76 3.185 1.64 3.305 1.64 3.305 1.54 3.705 1.54 3.705 1.18 3.185 1.18 3.185 0.9 3.005 0.9 3.005 0.66 3.125 0.66 3.125 0.78 3.305 0.78 3.305 1.06 4.285 1.06 ;
      POLYGON 3.785 0.52 2.785 0.52 2.785 0.78 2.705 0.78 2.705 0.9 2.665 0.9 2.665 1.28 2.825 1.28 2.825 1.82 2.705 1.82 2.705 1.4 2.545 1.4 2.545 0.78 2.585 0.78 2.585 0.66 2.665 0.66 2.665 0.4 3.785 0.4 ;
      POLYGON 3.585 1.42 3.065 1.42 3.065 2.06 2.465 2.06 2.465 1.64 1.865 1.64 1.865 1.82 1.745 1.82 1.745 1.38 1.585 1.38 1.585 0.66 1.705 0.66 1.705 1.26 1.865 1.26 1.865 1.52 2.585 1.52 2.585 1.94 2.945 1.94 2.945 1.16 2.785 1.16 2.785 1.04 3.065 1.04 3.065 1.3 3.585 1.3 ;
      POLYGON 1.465 1.675 1.155 1.675 1.155 1.77 0.915 1.77 0.915 1.675 0.415 1.675 0.415 1.27 0.535 1.27 0.535 1.555 1.345 1.555 1.345 0.765 1.135 0.765 1.135 0.645 1.465 0.645 ;
  END
END ADDHXL

MACRO DFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX4 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.49 2.175 1.61 ;
        RECT 1.935 1.315 2.14 1.61 ;
        RECT 2.02 0.63 2.14 1.61 ;
        RECT 1.23 1.315 2.14 1.435 ;
        RECT 1.18 1.175 1.38 1.315 ;
        RECT 0.975 1.49 1.35 1.61 ;
        RECT 1.23 1.175 1.35 1.61 ;
        RECT 1.18 0.63 1.3 1.315 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.88 0.93 9 1.24 ;
        RECT 8.77 0.83 8.92 1.145 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.11 0.855 1.38 ;
        RECT 0.495 1.11 0.855 1.36 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.755 1.16 6.535 1.28 ;
        RECT 6.415 1.04 6.535 1.28 ;
        RECT 5.755 0.36 5.875 1.28 ;
        RECT 4.615 0.36 5.875 0.48 ;
        RECT 3.505 0.73 4.735 0.85 ;
        RECT 4.615 0.36 4.735 0.85 ;
        RECT 3.695 0.73 3.815 1.1 ;
        RECT 3.505 0.36 3.625 0.85 ;
        RECT 2.71 0.36 3.625 0.48 ;
        RECT 2.71 0.36 2.83 1.12 ;
        RECT 2.68 0.595 2.83 0.855 ;
    END
  END RN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 8.94 -0.18 9.06 0.71 ;
        RECT 5.995 -0.18 6.115 0.68 ;
        RECT 3.835 0.49 4.075 0.61 ;
        RECT 3.835 -0.18 3.955 0.61 ;
        RECT 2.44 -0.18 2.56 0.68 ;
        RECT 1.6 -0.18 1.72 0.68 ;
        RECT 0.76 -0.18 0.88 0.87 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.04 1.6 9.16 2.79 ;
        RECT 7.36 2.29 7.6 2.79 ;
        RECT 5.86 2.25 6.1 2.79 ;
        RECT 4.215 1.94 4.335 2.79 ;
        RECT 3.315 2.23 3.435 2.79 ;
        RECT 2.475 2.23 2.595 2.79 ;
        RECT 1.455 1.97 1.695 2.09 ;
        RECT 1.455 1.97 1.575 2.79 ;
        RECT 0.495 1.97 0.735 2.09 ;
        RECT 0.495 1.97 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.58 1.84 9.46 1.84 9.46 1.72 9.36 1.72 9.36 1.48 8.76 1.48 8.76 2.2 8.05 2.2 8.05 1.93 6.655 1.93 6.655 1.89 5.095 1.89 5.095 1.33 4.655 1.33 4.655 1.21 5.095 1.21 5.095 1 5.275 1 5.275 0.88 5.395 0.88 5.395 1.12 5.215 1.12 5.215 1.77 6.775 1.77 6.775 1.81 8.05 1.81 8.05 1.32 7.635 1.32 7.635 1.16 7.515 1.16 7.515 1.04 7.755 1.04 7.755 1.2 8.17 1.2 8.17 2.08 8.64 2.08 8.64 1.385 8.53 1.385 8.53 1.1 8.65 1.1 8.65 1.265 8.76 1.265 8.76 1.36 9.36 1.36 9.36 0.47 9.48 0.47 9.48 1.6 9.58 1.6 ;
      POLYGON 8.52 1.96 8.4 1.96 8.4 1.625 8.29 1.625 8.29 0.92 6.235 0.92 6.235 1.04 5.995 1.04 5.995 0.8 7.735 0.8 7.735 0.54 7.855 0.54 7.855 0.8 8.41 0.8 8.41 1.505 8.52 1.505 ;
      POLYGON 7.93 1.69 7.81 1.69 7.81 1.65 7.135 1.65 7.135 1.69 6.895 1.69 6.895 1.53 7.81 1.53 7.81 1.44 7.93 1.44 ;
      POLYGON 7.92 2.17 6.415 2.17 6.415 2.13 5.74 2.13 5.74 2.23 5.315 2.23 5.315 2.25 5.075 2.25 5.075 2.23 4.56 2.23 4.56 1.82 4.095 1.82 4.095 2.11 1.99 2.11 1.99 1.85 0.375 1.85 0.375 1.91 0.255 1.91 0.255 2.03 0.135 2.03 0.135 1.73 0.255 1.73 0.255 0.69 0.52 0.69 0.52 0.81 0.375 0.81 0.375 1.73 2.11 1.73 2.11 1.99 3.975 1.99 3.975 1.7 4.68 1.7 4.68 2.11 5.62 2.11 5.62 2.01 6.535 2.01 6.535 2.05 7.92 2.05 ;
      POLYGON 7.355 1.41 6.775 1.41 6.775 1.52 5.635 1.52 5.635 1.65 5.335 1.65 5.335 1.53 5.515 1.53 5.515 0.72 5.375 0.72 5.375 0.6 5.635 0.6 5.635 1.4 6.655 1.4 6.655 1.29 7.235 1.29 7.235 1.11 7.355 1.11 ;
      POLYGON 5.195 0.72 4.975 0.72 4.975 1.09 4.535 1.09 4.535 1.45 4.92 1.45 4.92 1.57 4.975 1.57 4.975 1.99 4.855 1.99 4.855 1.69 4.8 1.69 4.8 1.57 4.415 1.57 4.415 1.09 4.055 1.09 4.055 1.34 3.335 1.34 3.335 1.1 3.455 1.1 3.455 1.22 3.935 1.22 3.935 0.97 4.855 0.97 4.855 0.6 5.195 0.6 ;
      POLYGON 4.295 1.58 3.855 1.58 3.855 1.87 3.615 1.87 3.615 1.72 3.735 1.72 3.735 1.58 2.955 1.58 2.955 1.87 2.835 1.87 2.835 1.36 2.275 1.36 2.275 1.11 2.395 1.11 2.395 1.24 2.955 1.24 2.955 1.46 3.095 1.46 3.095 0.6 3.375 0.6 3.375 0.72 3.215 0.72 3.215 1.46 4.175 1.46 4.175 1.34 4.295 1.34 ;
  END
END DFFRHQX4

MACRO NAND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1.055 0.815 1.485 ;
        RECT 0.65 0.885 0.8 1.3 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.355 1.06 0.51 1.515 ;
        RECT 0.355 1.04 0.475 1.515 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 1.025 1.175 1.265 ;
        RECT 0.94 0.885 1.115 1.145 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.485 1.605 1.605 1.845 ;
        RECT 0.63 1.605 1.605 1.725 ;
        RECT 1.23 1.465 1.415 1.725 ;
        RECT 1.295 0.68 1.415 1.725 ;
        RECT 0.495 1.635 0.75 1.755 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.195 -0.18 0.315 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 1.005 2.155 1.125 2.79 ;
        RECT 0.135 1.635 0.255 2.79 ;
    END
  END VDD
END NAND3XL

MACRO SEDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX4 0 0 ;
  SIZE 14.5 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.405 1.5 1.525 2.15 ;
        RECT 1.405 0.68 1.525 1.025 ;
        RECT 1.385 0.905 1.505 1.62 ;
        RECT 0.565 1.025 1.505 1.145 ;
        RECT 0.565 0.885 0.8 1.145 ;
        RECT 0.565 0.68 0.685 2.15 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.23 8.105 1.5 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.135 0.895 8.395 1.11 ;
        RECT 8.245 0.895 8.365 1.275 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.185 1.09 10.37 1.505 ;
        RECT 10.185 1.09 10.305 1.52 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.37 1.43 13.585 1.67 ;
        RECT 13.325 1.465 13.56 1.725 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.13 1.125 13.985 1.245 ;
        RECT 13.7 0.885 13.85 1.245 ;
        RECT 12.665 1.225 13.25 1.345 ;
        RECT 12.665 1.225 12.785 1.75 ;
    END
  END E
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.09 0.85 11.905 0.97 ;
        RECT 11.785 0.68 11.905 0.97 ;
        RECT 11.585 1.62 11.825 1.74 ;
        RECT 11.09 1.5 11.705 1.62 ;
        RECT 11.09 1.465 11.24 1.725 ;
        RECT 10.625 1.62 11.21 1.74 ;
        RECT 11.09 0.8 11.21 1.74 ;
        RECT 10.945 0.8 11.21 0.92 ;
        RECT 10.945 0.68 11.065 0.92 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 14.5 0.18 ;
        RECT 13.585 -0.18 13.705 0.765 ;
        RECT 12.205 -0.18 12.325 0.73 ;
        RECT 11.365 -0.18 11.485 0.73 ;
        RECT 10.525 -0.18 10.645 0.73 ;
        RECT 8.225 0.415 8.465 0.535 ;
        RECT 8.345 -0.18 8.465 0.535 ;
        RECT 6.79 -0.18 6.91 0.73 ;
        RECT 4.445 0.61 4.685 0.73 ;
        RECT 4.565 -0.18 4.685 0.73 ;
        RECT 2.725 -0.18 2.845 0.82 ;
        RECT 1.825 -0.18 1.945 0.73 ;
        RECT 0.985 -0.18 1.105 0.73 ;
        RECT 0.145 -0.18 0.265 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 14.5 2.79 ;
        RECT 13.625 2.085 13.745 2.79 ;
        RECT 12.065 2.1 12.305 2.22 ;
        RECT 12.065 2.1 12.185 2.79 ;
        RECT 11.105 2.1 11.345 2.22 ;
        RECT 11.105 2.1 11.225 2.79 ;
        RECT 10.145 2.1 10.385 2.22 ;
        RECT 10.145 2.1 10.265 2.79 ;
        RECT 8.235 1.86 8.355 2.79 ;
        RECT 6.645 1.88 6.765 2.79 ;
        RECT 6.525 1.88 6.765 2 ;
        RECT 4.625 1.81 4.745 2.79 ;
        RECT 4.505 1.81 4.745 1.93 ;
        RECT 2.725 2.02 2.845 2.79 ;
        RECT 1.825 1.63 1.945 2.79 ;
        RECT 0.985 1.5 1.105 2.79 ;
        RECT 0.145 1.5 0.265 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 14.225 2.09 14.105 2.09 14.105 1.965 13.065 1.965 13.065 1.53 13.185 1.53 13.185 1.845 14.105 1.845 14.105 1.005 14.005 1.005 14.005 0.525 14.125 0.525 14.125 0.885 14.225 0.885 ;
      POLYGON 13.065 0.97 12.545 0.97 12.545 1.87 12.945 1.87 12.945 2.11 12.825 2.11 12.825 1.99 12.425 1.99 12.425 1.98 9.295 1.98 9.295 1.38 9.585 1.38 9.585 0.86 9.505 0.86 9.505 0.6 9.625 0.6 9.625 0.74 9.705 0.74 9.705 1.5 9.415 1.5 9.415 1.86 12.425 1.86 12.425 0.85 12.945 0.85 12.945 0.525 13.065 0.525 ;
      POLYGON 10.785 1.24 10.665 1.24 10.665 1.09 10.55 1.09 10.55 0.97 10.285 0.97 10.285 0.56 9.84 0.56 9.84 0.48 8.9 0.48 8.9 0.775 7.985 0.775 7.985 0.48 7.33 0.48 7.33 0.8 7.485 0.8 7.485 1.77 7.365 1.77 7.365 0.92 7.21 0.92 7.21 0.36 8.105 0.36 8.105 0.655 8.78 0.655 8.78 0.36 9.96 0.36 9.96 0.44 10.405 0.44 10.405 0.85 10.67 0.85 10.67 0.97 10.785 0.97 ;
      POLYGON 10.165 0.92 9.945 0.92 9.945 1.74 9.665 1.74 9.665 1.62 9.825 1.62 9.825 0.8 10.045 0.8 10.045 0.68 10.165 0.68 ;
      POLYGON 9.465 1.26 8.965 1.26 8.965 1.6 8.725 1.6 8.725 1.48 8.845 1.48 8.845 1.14 9.345 1.14 9.345 0.98 9.465 0.98 ;
      POLYGON 9.205 1.02 8.635 1.02 8.635 1.36 8.605 1.36 8.605 1.8 9.055 1.8 9.055 1.92 8.485 1.92 8.485 1.74 8.115 1.74 8.115 2.25 6.885 2.25 6.885 1.76 5.745 1.76 5.745 1.87 5.625 1.87 5.625 1.61 5.805 1.61 5.805 0.86 5.745 0.86 5.745 0.62 5.865 0.62 5.865 0.74 5.925 0.74 5.925 1.64 7.005 1.64 7.005 2.13 7.995 2.13 7.995 1.62 8.485 1.62 8.485 1.24 8.515 1.24 8.515 0.9 9.085 0.9 9.085 0.6 9.205 0.6 ;
      POLYGON 7.875 2.01 7.125 2.01 7.125 1.2 6.325 1.2 6.325 1.08 7.245 1.08 7.245 1.89 7.605 1.89 7.605 0.99 7.745 0.99 7.745 0.6 7.865 0.6 7.865 1.11 7.725 1.11 7.725 1.74 7.875 1.74 ;
      POLYGON 6.43 0.92 6.205 0.92 6.205 1.4 6.285 1.4 6.285 1.52 6.045 1.52 6.045 1.4 6.085 1.4 6.085 0.8 6.31 0.8 6.31 0.68 6.045 0.68 6.045 0.5 5.625 0.5 5.625 1.37 5.685 1.37 5.685 1.49 5.445 1.49 5.445 1.37 5.505 1.37 5.505 0.5 4.925 0.5 4.925 0.97 4.205 0.97 4.205 0.5 3.365 0.5 3.365 1.18 3.385 1.18 3.385 1.42 3.245 1.42 3.245 0.38 3.765 0.38 3.765 0.36 4.005 0.36 4.005 0.38 4.325 0.38 4.325 0.85 4.805 0.85 4.805 0.38 5.005 0.38 5.005 0.36 5.245 0.36 5.245 0.38 6.165 0.38 6.165 0.56 6.43 0.56 ;
      POLYGON 6.405 2.2 5.395 2.2 5.395 2.11 4.865 2.11 4.865 1.69 4.385 1.69 4.385 2.11 3.745 2.11 3.745 2.05 3.245 2.05 3.245 2.25 3.005 2.25 3.005 1.9 2.365 1.9 2.365 2.15 2.245 2.15 2.245 1.75 2.205 1.75 2.205 1.36 1.625 1.36 1.625 1.24 2.205 1.24 2.205 0.8 2.305 0.8 2.305 0.68 2.425 0.68 2.425 0.92 2.325 0.92 2.325 1.63 2.365 1.63 2.365 1.78 3.125 1.78 3.125 1.93 3.865 1.93 3.865 1.99 4.265 1.99 4.265 1.57 4.985 1.57 4.985 1.99 5.515 1.99 5.515 2.08 6.405 2.08 ;
      POLYGON 5.385 0.8 5.265 0.8 5.265 1.63 5.325 1.63 5.325 1.87 5.205 1.87 5.205 1.75 5.145 1.75 5.145 1.21 4.225 1.21 4.225 1.09 5.145 1.09 5.145 0.68 5.385 0.68 ;
      POLYGON 4.905 1.45 4.105 1.45 4.105 1.87 3.985 1.87 3.985 1.21 3.965 1.21 3.965 0.62 4.085 0.62 4.085 1.09 4.105 1.09 4.105 1.33 4.905 1.33 ;
      POLYGON 3.745 1.81 3.505 1.81 3.505 1.66 3.005 1.66 3.005 1.47 2.445 1.47 2.445 1.35 3.125 1.35 3.125 1.54 3.505 1.54 3.505 0.8 3.485 0.8 3.485 0.68 3.725 0.68 3.725 0.8 3.625 0.8 3.625 1.69 3.745 1.69 ;
  END
END SEDFFX4

MACRO AND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.35 0.78 0.53 1.16 ;
        RECT 0.33 0.79 0.48 1.18 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.78 0.82 1.2 ;
        RECT 0.65 0.78 0.82 1.185 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.135 0.96 1.255 1.2 ;
        RECT 0.94 0.96 1.255 1.145 ;
        RECT 0.94 0.885 1.09 1.145 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.675 1.36 1.93 1.48 ;
        RECT 1.675 1.24 1.795 1.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 0.885 3.41 1.145 ;
        RECT 3.075 1.32 3.195 2.21 ;
        RECT 3.055 0.68 3.175 1.44 ;
        RECT 2.235 1.32 3.195 1.44 ;
        RECT 2.095 0.73 3.175 0.85 ;
        RECT 2.815 0.68 3.175 0.85 ;
        RECT 2.235 1.32 2.355 2.21 ;
        RECT 1.975 0.68 2.215 0.8 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.295 -0.18 3.415 0.67 ;
        RECT 2.395 0.49 2.635 0.61 ;
        RECT 2.395 -0.18 2.515 0.61 ;
        RECT 1.615 -0.18 1.735 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.495 1.56 3.615 2.79 ;
        RECT 2.655 1.56 2.775 2.79 ;
        RECT 1.815 1.845 1.935 2.79 ;
        RECT 0.975 1.56 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.935 1.14 2.695 1.14 2.695 1.12 2.475 1.12 2.475 1.14 2.235 1.14 2.235 1.12 1.495 1.12 1.495 1.32 1.515 1.32 1.515 2.21 1.395 2.21 1.395 1.44 0.675 1.44 0.675 2.21 0.555 2.21 0.555 1.32 1.375 1.32 1.375 0.66 0.16 0.66 0.16 0.54 1.495 0.54 1.495 1 2.815 1 2.815 1.02 2.935 1.02 ;
  END
END AND4X4

MACRO OR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X8 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.95 2.135 1.13 ;
        RECT 1.755 0.94 2.015 1.13 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.255 1.25 2.595 1.37 ;
        RECT 2.475 0.94 2.595 1.37 ;
        RECT 2.335 0.94 2.595 1.09 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.49 2.975 1.61 ;
        RECT 2.855 1.24 2.975 1.61 ;
        RECT 0.68 1.28 1.075 1.61 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 1.52 3.465 1.67 ;
        RECT 0.41 1.73 3.335 1.85 ;
        RECT 3.215 1.22 3.335 1.85 ;
        RECT 3.205 1.52 3.335 1.85 ;
        RECT 0.41 1.22 0.53 1.85 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.335 0.715 6.695 0.835 ;
        RECT 6.415 1.23 6.535 2.21 ;
        RECT 4.055 0.765 6.455 0.885 ;
        RECT 5.695 1.23 6.535 1.35 ;
        RECT 5.695 0.765 6.02 1.35 ;
        RECT 3.895 1.275 5.815 1.395 ;
        RECT 5.675 0.645 5.795 0.885 ;
        RECT 5.575 1.275 5.695 2.21 ;
        RECT 4.775 0.715 5.015 0.885 ;
        RECT 4.735 1.275 4.855 2.21 ;
        RECT 3.935 0.715 4.175 0.835 ;
        RECT 3.895 1.275 4.015 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.095 -0.18 6.215 0.645 ;
        RECT 5.255 -0.18 5.375 0.645 ;
        RECT 4.415 -0.18 4.535 0.645 ;
        RECT 3.515 0.46 3.755 0.58 ;
        RECT 3.515 -0.18 3.635 0.58 ;
        RECT 2.675 0.46 2.915 0.58 ;
        RECT 2.675 -0.18 2.795 0.58 ;
        RECT 1.835 0.46 2.075 0.58 ;
        RECT 1.835 -0.18 1.955 0.58 ;
        RECT 0.995 0.46 1.235 0.58 ;
        RECT 0.995 -0.18 1.115 0.58 ;
        RECT 0.215 -0.18 0.335 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 5.995 1.47 6.115 2.79 ;
        RECT 5.155 1.515 5.275 2.79 ;
        RECT 4.315 1.515 4.435 2.79 ;
        RECT 3.355 2.21 3.595 2.79 ;
        RECT 0.415 1.97 0.535 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.575 1.155 3.705 1.155 3.705 2.09 2.175 2.09 2.175 2.15 1.935 2.15 1.935 1.97 3.585 1.97 3.585 0.82 0.695 0.82 0.695 0.77 0.575 0.77 0.575 0.65 0.815 0.65 0.815 0.7 1.415 0.7 1.415 0.65 1.655 0.65 1.655 0.7 2.255 0.7 2.255 0.65 2.495 0.65 2.495 0.7 3.095 0.7 3.095 0.65 3.335 0.65 3.335 0.7 3.705 0.7 3.705 1.035 5.575 1.035 ;
  END
END OR4X8

MACRO DFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX1 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.635 0.85 4.755 1.15 ;
        RECT 4.235 0.85 4.755 0.97 ;
        RECT 4.235 0.36 4.355 0.97 ;
        RECT 2.39 0.36 4.355 0.48 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.39 0.36 2.51 1.34 ;
        RECT 1.97 1.22 2.51 1.34 ;
        RECT 1.85 1.26 2.09 1.38 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.975 1.12 7.235 1.39 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 1.165 7.815 1.38 ;
        RECT 7.435 1.12 7.675 1.31 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.64 0.54 1.99 ;
        RECT 0.07 1.175 0.54 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.295 -0.18 7.415 0.74 ;
        RECT 5.715 0.46 5.955 0.58 ;
        RECT 5.715 -0.18 5.835 0.58 ;
        RECT 4.475 0.61 4.715 0.73 ;
        RECT 4.475 -0.18 4.595 0.73 ;
        RECT 1.65 -0.18 1.77 0.68 ;
        RECT 0.84 -0.18 0.96 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.095 1.75 7.215 2.79 ;
        RECT 5.735 1.68 5.855 2.79 ;
        RECT 4.655 2.23 4.895 2.79 ;
        RECT 2.43 1.98 2.67 2.15 ;
        RECT 2.43 1.98 2.55 2.79 ;
        RECT 1.65 1.74 1.77 2.79 ;
        RECT 0.84 1.34 0.96 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.835 0.88 7.655 0.88 7.655 1 6.855 1 6.855 1.51 7.505 1.51 7.505 1.66 7.635 1.66 7.635 1.9 7.515 1.9 7.515 1.78 7.385 1.78 7.385 1.63 6.975 1.63 6.975 2.21 6.395 2.21 6.395 2.25 6.155 2.25 6.155 2.13 6.205 2.13 6.205 1.56 5.615 1.56 5.615 2.21 5.015 2.21 5.015 2.11 4.335 2.11 4.335 1.99 5.135 1.99 5.135 2.09 5.495 2.09 5.495 1.44 6.325 1.44 6.325 2.09 6.735 2.09 6.735 0.88 7.535 0.88 7.535 0.76 7.715 0.76 7.715 0.5 7.835 0.5 ;
      POLYGON 6.635 0.76 6.615 0.76 6.615 1.32 6.575 1.32 6.575 1.97 6.455 1.97 6.455 1.32 5.475 1.32 5.475 1.19 5.715 1.19 5.715 1.2 6.495 1.2 6.495 0.64 6.515 0.64 6.515 0.5 6.635 0.5 ;
      POLYGON 6.375 1.08 6.255 1.08 6.255 0.83 5.475 0.83 5.475 0.53 4.995 0.53 4.995 1.39 4.295 1.39 4.295 1.51 4.415 1.51 4.415 1.63 4.175 1.63 4.175 1.21 3.98 1.21 3.98 0.73 3.875 0.73 3.875 0.61 4.115 0.61 4.115 0.73 4.1 0.73 4.1 1.09 4.295 1.09 4.295 1.27 4.875 1.27 4.875 0.41 5.595 0.41 5.595 0.71 6.375 0.71 ;
      POLYGON 6.075 1.07 5.355 1.07 5.355 1.45 5.375 1.45 5.375 1.97 5.255 1.97 5.255 1.87 3.92 1.87 3.92 2.21 3.8 2.21 3.8 1.45 3.74 1.45 3.74 0.97 3.05 0.97 3.05 0.6 3.29 0.6 3.29 0.85 3.86 0.85 3.86 1.33 3.92 1.33 3.92 1.75 5.255 1.75 5.255 1.57 5.235 1.57 5.235 0.77 5.115 0.77 5.115 0.65 5.355 0.65 5.355 0.95 6.075 0.95 ;
      POLYGON 3.62 1.34 2.9 1.34 2.9 1.1 3.02 1.1 3.02 1.22 3.62 1.22 ;
      POLYGON 3.5 2.21 3.38 2.21 3.38 1.58 2.78 1.58 2.78 1.62 1.51 1.62 1.51 1.37 1.63 1.37 1.63 1.5 2.66 1.5 2.66 0.72 2.63 0.72 2.63 0.6 2.87 0.6 2.87 0.72 2.78 0.72 2.78 1.46 3.5 1.46 ;
      POLYGON 3.08 2.21 2.96 2.21 2.96 1.86 2.19 1.86 2.19 2.21 2.07 2.21 2.07 1.74 2.96 1.74 2.96 1.7 3.08 1.7 ;
      POLYGON 2.27 1.1 1.35 1.1 1.35 2.21 1.23 2.21 1.23 1.1 0.8 1.1 0.8 1.22 0.68 1.22 0.68 0.98 1.23 0.98 1.23 0.54 1.35 0.54 1.35 0.98 2.15 0.98 2.15 0.86 2.27 0.86 ;
  END
END DFFSHQX1

MACRO SDFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX1 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.43 4.025 1.55 ;
        RECT 2.845 1.75 3.905 1.87 ;
        RECT 3.785 1.43 3.905 1.87 ;
        RECT 2.845 1.75 2.965 2.01 ;
        RECT 2.315 1.89 2.965 2.01 ;
        RECT 1.575 1.99 2.435 2.11 ;
        RECT 1.575 1.35 1.73 1.59 ;
        RECT 1.575 1.35 1.695 2.11 ;
        RECT 1.52 1.465 1.695 1.725 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.245 1.23 7.61 1.39 ;
        RECT 7.245 1.23 7.605 1.425 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.41 0.94 7.825 1.11 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.005 1.2 9.265 1.43 ;
        RECT 9.105 1.2 9.225 1.61 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.715 0.96 9.835 1.2 ;
        RECT 9.64 0.885 9.79 1.145 ;
        RECT 8.485 0.96 9.835 1.08 ;
        RECT 8.485 0.96 8.725 1.09 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2696 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.675 1.22 1.09 1.34 ;
        RECT 0.675 0.72 0.915 0.84 ;
        RECT 0.675 0.72 0.795 1.46 ;
        RECT 0.605 1.34 0.725 1.58 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 9.995 -0.18 10.115 0.765 ;
        RECT 9.105 -0.18 9.225 0.6 ;
        RECT 7.625 0.46 7.865 0.58 ;
        RECT 7.745 -0.18 7.865 0.58 ;
        RECT 6.425 -0.18 6.665 0.34 ;
        RECT 4.825 -0.18 4.945 0.75 ;
        RECT 3.645 -0.18 3.765 0.65 ;
        RECT 1.53 0.5 1.77 0.62 ;
        RECT 1.53 -0.18 1.65 0.62 ;
        RECT 0.075 0.53 0.315 0.65 ;
        RECT 0.075 -0.18 0.195 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 10.055 1.98 10.175 2.79 ;
        RECT 9.265 1.97 9.385 2.79 ;
        RECT 7.685 1.56 7.805 2.79 ;
        RECT 6.755 1.46 6.875 2.79 ;
        RECT 4.595 2.23 4.835 2.79 ;
        RECT 3.635 2.23 3.875 2.79 ;
        RECT 2.295 2.23 2.535 2.79 ;
        RECT 1.335 2.23 1.575 2.79 ;
        RECT 0.185 1.34 0.305 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.755 0.705 9.52 0.705 9.52 0.84 8.365 0.84 8.365 1.21 8.885 1.21 8.885 1.73 9.345 1.73 9.345 1.55 9.515 1.55 9.515 1.52 9.755 1.52 9.755 1.67 9.465 1.67 9.465 1.85 8.765 1.85 8.765 1.33 8.185 1.33 8.185 0.94 8.245 0.94 8.245 0.72 9.4 0.72 9.4 0.585 9.755 0.585 ;
      POLYGON 8.745 2.21 8.625 2.21 8.625 2.09 8.525 2.09 8.525 1.57 7.945 1.57 7.945 0.82 7.385 0.82 7.385 0.53 6.905 0.53 6.905 0.58 6.155 0.58 6.155 1.79 6.175 1.79 6.175 2.01 5.935 2.01 5.935 1.79 6.035 1.79 6.035 0.81 5.945 0.81 5.945 0.46 6.785 0.46 6.785 0.41 7.505 0.41 7.505 0.7 8 0.7 8 0.48 8.505 0.48 8.505 0.6 8.12 0.6 8.12 0.82 8.065 0.82 8.065 1.45 8.645 1.45 8.645 1.97 8.745 1.97 ;
      POLYGON 7.325 1.8 7.205 1.8 7.205 1.665 7.005 1.665 7.005 1.19 6.555 1.19 6.555 1.07 7.005 1.07 7.005 0.7 7.025 0.7 7.025 0.65 7.265 0.65 7.265 0.82 7.125 0.82 7.125 1.545 7.325 1.545 ;
      POLYGON 6.515 0.86 6.435 0.86 6.435 1.34 6.455 1.34 6.455 2.25 5.165 2.25 5.165 2.11 3.205 2.11 3.205 2.25 2.805 2.25 2.805 2.13 3.085 2.13 3.085 1.99 5.285 1.99 5.285 2.13 5.695 2.13 5.695 1.37 5.815 1.37 5.815 2.13 6.335 2.13 6.335 1.46 6.315 1.46 6.315 0.86 6.275 0.86 6.275 0.74 6.515 0.74 ;
      POLYGON 5.915 1.17 5.795 1.17 5.795 1.05 5.705 1.05 5.705 0.49 5.335 0.49 5.335 1.57 5.215 1.57 5.215 0.99 4.585 0.99 4.585 0.48 4.175 0.48 4.175 0.89 3.49 0.89 3.49 0.99 3.37 0.99 3.37 0.48 2.45 0.48 2.45 0.88 2.55 0.88 2.55 1.12 2.33 1.12 2.33 0.36 3.49 0.36 3.49 0.77 4.055 0.77 4.055 0.36 4.705 0.36 4.705 0.87 5.215 0.87 5.215 0.37 5.825 0.37 5.825 0.93 5.915 0.93 ;
      POLYGON 5.585 0.85 5.575 0.85 5.575 1.81 5.535 1.81 5.535 2.01 5.415 2.01 5.415 1.81 4.475 1.81 4.475 1.59 4.435 1.59 4.435 1.35 4.555 1.35 4.555 1.47 4.595 1.47 4.595 1.69 5.455 1.69 5.455 0.73 5.465 0.73 5.465 0.61 5.585 0.61 ;
      POLYGON 5.055 1.23 4.315 1.23 4.315 1.75 4.355 1.75 4.355 1.87 4.115 1.87 4.115 1.75 4.195 1.75 4.195 1.23 3.565 1.23 3.565 1.63 3.445 1.63 3.445 1.23 3.13 1.23 3.13 0.72 2.99 0.72 2.99 0.6 3.25 0.6 3.25 1.11 4.345 1.11 4.345 0.6 4.465 0.6 4.465 1.11 5.055 1.11 ;
      POLYGON 3.145 1.63 3.025 1.63 3.025 1.47 2.89 1.47 2.89 1.36 1.85 1.36 1.85 1.19 1.45 1.19 1.45 1.07 1.97 1.07 1.97 1.24 2.67 1.24 2.67 0.72 2.57 0.72 2.57 0.6 2.81 0.6 2.81 0.72 2.79 0.72 2.79 1.24 3.01 1.24 3.01 1.35 3.145 1.35 ;
      POLYGON 2.725 1.77 2.055 1.77 2.055 1.87 1.815 1.87 1.815 1.75 1.935 1.75 1.935 1.65 2.605 1.65 2.605 1.48 2.725 1.48 ;
      POLYGON 2.21 1.1 2.09 1.1 2.09 0.86 1.33 0.86 1.33 1.675 1.035 1.675 1.035 2.21 0.915 2.21 0.915 1.555 1.21 1.555 1.21 0.86 1.035 0.86 1.035 0.6 0.555 0.6 0.555 1.22 0.435 1.22 0.435 0.48 1.155 0.48 1.155 0.54 1.29 0.54 1.29 0.66 1.33 0.66 1.33 0.74 2.21 0.74 ;
  END
END SDFFSHQX1

MACRO SDFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX4 0 0 ;
  SIZE 12.18 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.33 1.515 2.08 ;
        RECT 1.395 0.63 1.515 0.97 ;
        RECT 1.375 0.85 1.495 1.45 ;
        RECT 0.555 0.97 1.495 1.09 ;
        RECT 0.555 0.885 0.8 1.145 ;
        RECT 0.555 0.63 0.675 2.08 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.205 1.4 5.445 1.52 ;
        RECT 5.205 1.4 5.325 1.76 ;
        RECT 4.615 1.72 5.265 1.84 ;
        RECT 5.145 1.64 5.325 1.76 ;
        RECT 4.085 1.89 4.735 2.01 ;
        RECT 4.615 1.72 4.735 2.01 ;
        RECT 4.085 1.7 4.205 2.01 ;
        RECT 3.375 1.7 4.205 1.82 ;
        RECT 2.71 1.99 3.495 2.11 ;
        RECT 3.375 1.7 3.495 2.11 ;
        RECT 2.675 1.17 2.915 1.29 ;
        RECT 2.71 1.17 2.83 2.11 ;
        RECT 2.68 1.465 2.83 1.725 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.715 1.21 8.975 1.45 ;
        RECT 8.645 1.115 8.885 1.33 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.515 0.94 9.635 1.18 ;
        RECT 9.005 0.94 9.635 1.06 ;
        RECT 9.005 0.94 9.265 1.09 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.035 1.22 11.31 1.415 ;
        RECT 11.035 1.22 11.165 1.555 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.355 0.98 11.91 1.1 ;
        RECT 11.67 0.885 11.82 1.145 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.18 0.18 ;
        RECT 11.925 -0.18 12.045 0.765 ;
        RECT 10.975 -0.18 11.095 0.62 ;
        RECT 9.495 0.46 9.735 0.58 ;
        RECT 9.615 -0.18 9.735 0.58 ;
        RECT 8.295 -0.18 8.535 0.32 ;
        RECT 6.305 -0.18 6.425 0.68 ;
        RECT 5.125 -0.18 5.245 0.72 ;
        RECT 2.655 0.45 2.895 0.57 ;
        RECT 2.655 -0.18 2.775 0.57 ;
        RECT 1.815 -0.18 1.935 0.68 ;
        RECT 0.975 -0.18 1.095 0.68 ;
        RECT 0.135 -0.18 0.255 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.18 2.79 ;
        RECT 11.925 1.475 12.045 2.79 ;
        RECT 11.195 1.915 11.315 2.79 ;
        RECT 9.635 1.56 9.755 2.79 ;
        RECT 8.165 1.46 8.285 2.79 ;
        RECT 6.055 2.2 6.295 2.79 ;
        RECT 5.095 2.2 5.335 2.79 ;
        RECT 3.615 1.94 3.735 2.79 ;
        RECT 2.715 2.23 2.835 2.79 ;
        RECT 1.875 2.23 1.995 2.79 ;
        RECT 0.975 1.43 1.095 2.79 ;
        RECT 0.135 1.43 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.685 0.705 11.55 0.705 11.55 0.86 10.235 0.86 10.235 1.3 10.875 1.3 10.875 1.42 10.235 1.42 10.235 1.675 11.445 1.675 11.445 1.535 11.685 1.535 11.685 1.655 11.565 1.655 11.565 1.795 10.115 1.795 10.115 1.09 9.995 1.09 9.995 0.97 10.115 0.97 10.115 0.74 11.43 0.74 11.43 0.585 11.685 0.585 ;
      POLYGON 10.675 2.21 10.555 2.21 10.555 2.035 9.875 2.035 9.875 1.44 9.755 1.44 9.755 0.82 9.255 0.82 9.255 0.53 8.775 0.53 8.775 0.56 7.605 0.56 7.605 1.84 7.535 1.84 7.535 2.01 7.295 2.01 7.295 1.72 7.485 1.72 7.485 0.44 8.655 0.44 8.655 0.41 9.375 0.41 9.375 0.7 9.87 0.7 9.87 0.5 10.375 0.5 10.375 0.62 9.99 0.62 9.99 0.82 9.875 0.82 9.875 1.32 9.995 1.32 9.995 1.915 10.675 1.915 ;
      POLYGON 9.135 0.8 8.525 0.8 8.525 1.57 9.135 1.57 9.135 1.81 9.015 1.81 9.015 1.69 8.405 1.69 8.405 1.12 7.965 1.12 7.965 1 8.405 1 8.405 0.68 8.895 0.68 8.895 0.65 9.135 0.65 ;
      POLYGON 8.055 0.8 7.845 0.8 7.845 1.34 7.865 1.34 7.865 2.25 6.445 2.25 6.445 2.08 4.975 2.08 4.975 2.25 4.125 2.25 4.125 2.13 4.855 2.13 4.855 1.96 6.565 1.96 6.565 2.13 7.055 2.13 7.055 1.34 7.175 1.34 7.175 2.13 7.745 2.13 7.745 1.46 7.725 1.46 7.725 0.68 8.055 0.68 ;
      POLYGON 7.365 1.1 7.245 1.1 7.245 0.48 6.695 0.48 6.695 1.28 6.455 1.28 6.455 1.16 6.575 1.16 6.575 0.92 6.065 0.92 6.065 0.52 5.485 0.52 5.485 0.96 4.705 0.96 4.705 0.48 3.635 0.48 3.635 0.94 3.795 0.94 3.795 1.06 3.515 1.06 3.515 0.36 4.825 0.36 4.825 0.84 5.365 0.84 5.365 0.4 6.185 0.4 6.185 0.8 6.575 0.8 6.575 0.36 7.365 0.36 ;
      POLYGON 7.125 0.72 6.935 0.72 6.935 2.01 6.815 2.01 6.815 1.52 5.955 1.52 5.955 1.56 5.835 1.56 5.835 1.32 5.955 1.32 5.955 1.4 6.815 1.4 6.815 0.6 7.125 0.6 ;
      POLYGON 6.335 1.2 5.715 1.2 5.715 1.72 5.815 1.72 5.815 1.84 5.575 1.84 5.575 1.72 5.595 1.72 5.595 1.2 4.885 1.2 4.885 1.6 4.765 1.6 4.765 1.2 4.465 1.2 4.465 0.72 4.175 0.72 4.175 0.6 4.585 0.6 4.585 1.08 5.825 1.08 5.825 0.76 5.705 0.76 5.705 0.64 5.945 0.64 5.945 1.08 6.335 1.08 ;
      POLYGON 4.465 1.77 4.345 1.77 4.345 1.44 4.225 1.44 4.225 1.34 3.035 1.34 3.035 1.05 2.315 1.05 2.315 0.93 3.155 0.93 3.155 1.22 3.915 1.22 3.915 0.72 3.755 0.72 3.755 0.6 4.035 0.6 4.035 1.22 4.345 1.22 4.345 1.32 4.465 1.32 ;
      POLYGON 4.105 1.58 3.255 1.58 3.255 1.87 3.135 1.87 3.135 1.46 4.105 1.46 ;
      POLYGON 3.395 1.1 3.275 1.1 3.275 0.81 2.195 0.81 2.195 1.43 2.355 1.43 2.355 1.95 2.235 1.95 2.235 1.55 2.075 1.55 2.075 1.21 1.615 1.21 1.615 1.09 2.075 1.09 2.075 0.66 2.235 0.66 2.235 0.54 2.355 0.54 2.355 0.69 3.395 0.69 ;
  END
END SDFFSHQX4

MACRO TLATNTSCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX2 0 0 ;
  SIZE 6.67 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.325 0.82 0.565 1.22 ;
        RECT 0.305 0.82 0.565 1.09 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.76 1.09 1.175 ;
        RECT 0.925 0.81 1.045 1.245 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.76 1.38 1.22 ;
        RECT 1.245 0.76 1.365 1.245 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.995 0.59 6.115 0.83 ;
        RECT 5.87 0.71 6.02 1.145 ;
        RECT 5.865 1.145 5.99 1.265 ;
        RECT 5.865 1.145 5.985 1.99 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.67 0.18 ;
        RECT 6.415 -0.18 6.535 0.64 ;
        RECT 5.515 -0.18 5.635 0.53 ;
        RECT 4.655 -0.18 4.775 0.4 ;
        RECT 3.185 0.7 3.425 0.82 ;
        RECT 3.225 -0.18 3.345 0.82 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.67 2.79 ;
        RECT 6.285 1.34 6.405 2.79 ;
        RECT 5.445 1.36 5.565 2.79 ;
        RECT 4.605 1.48 4.725 2.79 ;
        RECT 3.025 2.14 3.265 2.26 ;
        RECT 3.025 2.14 3.145 2.79 ;
        RECT 0.925 1.605 1.045 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.745 1.18 5.185 1.18 5.185 1.44 5.145 1.44 5.145 1.6 5.025 1.6 5.025 1.32 5.065 1.32 5.065 1.06 5.305 1.06 5.305 0.86 5.185 0.86 5.185 0.74 5.425 0.74 5.425 1.06 5.745 1.06 ;
      POLYGON 5.265 0.52 5.065 0.52 5.065 0.64 4.415 0.64 4.415 0.56 3.945 0.56 3.945 0.76 3.905 0.76 3.905 1.3 2.945 1.3 2.945 1.66 3.745 1.66 3.745 1.89 3.865 1.89 3.865 2.01 3.625 2.01 3.625 1.78 2.825 1.78 2.825 1.3 2.685 1.3 2.685 1.18 3.785 1.18 3.785 0.64 3.825 0.64 3.825 0.44 4.535 0.44 4.535 0.52 4.945 0.52 4.945 0.4 5.265 0.4 ;
      POLYGON 4.945 1.2 4.295 1.2 4.295 1.42 4.305 1.42 4.305 1.66 4.185 1.66 4.185 1.54 3.065 1.54 3.065 1.42 4.175 1.42 4.175 0.68 4.295 0.68 4.295 1.08 4.945 1.08 ;
      POLYGON 4.465 2.25 3.385 2.25 3.385 2.02 2.505 2.02 2.505 2.07 2.385 2.07 2.385 1.95 2.205 1.95 2.205 0.64 2.325 0.64 2.325 1.83 2.505 1.83 2.505 1.9 3.505 1.9 3.505 2.13 4.345 2.13 4.345 1.82 4.465 1.82 ;
      POLYGON 3.705 0.48 3.665 0.48 3.665 1.06 2.945 1.06 2.945 0.52 2.565 0.52 2.565 1.57 2.705 1.57 2.705 1.69 2.445 1.69 2.445 0.52 1.62 0.52 1.62 1.605 1.525 1.605 1.525 1.725 1.405 1.725 1.405 1.485 1.5 1.485 1.5 0.64 1.395 0.64 1.395 0.4 1.985 0.4 1.985 0.36 2.225 0.36 2.225 0.4 3.065 0.4 3.065 0.94 3.545 0.94 3.545 0.48 3.465 0.48 3.465 0.36 3.705 0.36 ;
      POLYGON 2.085 2.07 1.965 2.07 1.965 1.965 1.165 1.965 1.165 1.485 0.405 1.485 0.405 1.725 0.285 1.725 0.285 1.365 0.685 1.365 0.685 0.7 0.555 0.7 0.555 0.4 0.675 0.4 0.675 0.58 0.805 0.58 0.805 1.365 1.285 1.365 1.285 1.845 1.965 1.845 1.965 0.88 1.785 0.88 1.785 0.64 1.905 0.64 1.905 0.76 2.085 0.76 ;
  END
END TLATNTSCAX2

MACRO XNOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 1.21 2.235 1.345 ;
        RECT 1.755 1.21 2.015 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.755 0.9 3.875 1.14 ;
        RECT 3.275 0.97 3.875 1.09 ;
        RECT 3.495 0.94 3.875 1.09 ;
        RECT 2.595 1.21 3.395 1.33 ;
        RECT 3.275 0.97 3.395 1.33 ;
        RECT 3.095 1.21 3.335 1.41 ;
        RECT 2.595 0.93 2.715 1.33 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 1.74 1.575 2.21 ;
        RECT 1.395 0.61 1.515 0.85 ;
        RECT 1.275 1.74 1.575 1.86 ;
        RECT 1.275 1.32 1.395 1.86 ;
        RECT 1.215 0.73 1.515 0.85 ;
        RECT 0.65 0.84 1.335 0.96 ;
        RECT 0.65 1.32 1.395 1.44 ;
        RECT 0.65 1.175 0.8 1.44 ;
        RECT 0.65 0.73 0.77 1.56 ;
        RECT 0.615 1.44 0.735 2.21 ;
        RECT 0.495 0.73 0.77 0.85 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.475 0.42 3.715 0.54 ;
        RECT 3.475 -0.18 3.595 0.54 ;
        RECT 1.755 0.54 1.995 0.66 ;
        RECT 1.755 -0.18 1.875 0.66 ;
        RECT 0.975 -0.18 1.095 0.72 ;
        RECT 0.135 -0.18 0.255 0.72 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.655 1.77 3.775 2.79 ;
        RECT 1.815 2.01 2.055 2.15 ;
        RECT 1.815 2.01 1.935 2.79 ;
        RECT 1.035 1.56 1.155 2.79 ;
        RECT 0.195 1.56 0.315 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.255 1.95 4.015 1.95 4.015 0.78 3.42 0.78 3.42 0.82 3.155 0.82 3.155 1.09 2.915 1.09 2.915 0.97 3.035 0.97 3.035 0.7 3.3 0.7 3.3 0.66 4.015 0.66 4.015 0.56 4.135 0.56 4.135 1.83 4.255 1.83 ;
      POLYGON 3.635 1.65 2.775 1.65 2.775 2.01 2.535 2.01 2.535 1.65 2.355 1.65 2.355 0.65 2.595 0.65 2.595 0.77 2.475 0.77 2.475 1.53 3.515 1.53 3.515 1.24 3.635 1.24 ;
      POLYGON 3.135 2.25 2.22 2.25 2.22 1.89 1.955 1.89 1.955 1.62 1.515 1.62 1.515 1.2 1.255 1.2 1.255 1.08 1.515 1.08 1.515 0.97 2.115 0.97 2.115 0.41 2.895 0.41 2.895 0.46 3.015 0.46 3.015 0.58 2.775 0.58 2.775 0.53 2.235 0.53 2.235 1.09 1.635 1.09 1.635 1.5 2.075 1.5 2.075 1.77 2.34 1.77 2.34 2.13 3.015 2.13 3.015 1.77 3.135 1.77 ;
  END
END XNOR2X4

MACRO DFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX2 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.05 0.51 1.52 ;
        RECT 0.39 1.02 0.51 1.52 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.08 0.835 1.51 ;
        RECT 0.65 1.145 0.8 1.56 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 1.465 5.73 1.725 ;
        RECT 5.58 1.13 5.7 1.725 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.61 1.175 7.76 1.435 ;
        RECT 7.635 1.175 7.755 2.16 ;
        RECT 7.61 0.74 7.73 1.435 ;
        RECT 7.455 0.74 7.73 0.86 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.415 0.74 8.655 0.86 ;
        RECT 8.48 1.175 8.63 1.435 ;
        RECT 8.48 0.74 8.6 1.435 ;
        RECT 8.475 1.295 8.595 2.16 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.895 -0.18 9.135 0.32 ;
        RECT 7.935 -0.18 8.175 0.38 ;
        RECT 6.975 -0.18 7.215 0.38 ;
        RECT 5.405 0.41 5.645 0.53 ;
        RECT 5.525 -0.18 5.645 0.53 ;
        RECT 1.615 -0.18 1.855 0.32 ;
        RECT 0.615 -0.18 0.735 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.895 1.51 9.015 2.79 ;
        RECT 8.055 1.51 8.175 2.79 ;
        RECT 7.215 1.64 7.335 2.79 ;
        RECT 6.405 2.09 6.525 2.79 ;
        RECT 5.665 2.09 5.785 2.79 ;
        RECT 4.64 2.29 4.88 2.79 ;
        RECT 1.955 2.2 2.075 2.79 ;
        RECT 0.655 1.68 0.775 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.495 0.86 9.435 0.86 9.435 1.75 9.315 1.75 9.315 1.29 8.75 1.29 8.75 1.17 9.315 1.17 9.315 0.86 9.255 0.86 9.255 0.74 9.495 0.74 ;
      POLYGON 9.415 0.62 8 0.62 8 1.24 7.88 1.24 7.88 0.62 7.335 0.62 7.335 1.06 7.455 1.06 7.455 1.18 7.115 1.18 7.115 1.52 6.975 1.52 6.975 2.1 6.735 2.1 6.735 1.7 6.855 1.7 6.855 1.4 6.995 1.4 6.995 1.04 6.155 1.04 6.155 0.92 6.555 0.92 6.555 0.68 6.675 0.68 6.675 0.92 7.215 0.92 7.215 0.5 9.295 0.5 9.295 0.36 9.415 0.36 ;
      POLYGON 6.875 1.28 5.915 1.28 5.915 1.01 5.46 1.01 5.46 1.24 4.625 1.24 4.625 1.12 5.34 1.12 5.34 0.89 6.035 0.89 6.035 1.16 6.875 1.16 ;
      POLYGON 6.345 0.72 6.225 0.72 6.225 0.77 5.065 0.77 5.065 0.48 4.585 0.48 4.585 0.6 4.265 0.6 4.265 0.82 4.025 0.82 4.025 0.7 4.145 0.7 4.145 0.48 4.465 0.48 4.465 0.36 5.185 0.36 5.185 0.65 6.105 0.65 6.105 0.6 6.345 0.6 ;
      POLYGON 6.145 1.965 5.34 1.965 5.34 1.93 4.265 1.93 4.265 1.82 4.145 1.82 4.145 1.7 4.385 1.7 4.385 1.81 5.46 1.81 5.46 1.845 6.025 1.845 6.025 1.57 6.145 1.57 ;
      POLYGON 5.305 1.69 5.185 1.69 5.185 1.57 4.505 1.57 4.505 1.58 4.025 1.58 4.025 1.98 2.435 1.98 2.435 1.4 2.195 1.4 2.195 1.28 2.555 1.28 2.555 1.86 3.165 1.86 3.165 1.74 3.125 1.74 3.125 0.76 3.185 0.76 3.185 0.64 3.305 0.64 3.305 0.88 3.245 0.88 3.245 1.62 3.285 1.62 3.285 1.86 3.905 1.86 3.905 1.46 4.385 1.46 4.385 0.72 4.705 0.72 4.705 0.6 4.945 0.6 4.945 0.72 4.825 0.72 4.825 0.84 4.505 0.84 4.505 1.45 5.305 1.45 ;
      POLYGON 5.22 2.17 4.305 2.17 4.305 2.22 2.195 2.22 2.195 2.04 1.415 2.04 1.415 1.8 1.335 1.8 1.335 0.84 1.215 0.84 1.215 0.72 1.455 0.72 1.455 1.68 1.535 1.68 1.535 1.92 2.315 1.92 2.315 2.1 4.185 2.1 4.185 2.05 5.22 2.05 ;
      POLYGON 4.265 1.34 3.785 1.34 3.785 1.7 3.525 1.7 3.525 1.58 3.665 1.58 3.665 0.64 3.785 0.64 3.785 1.22 4.265 1.22 ;
      POLYGON 4.005 0.48 3.885 0.48 3.885 0.5 3.545 0.5 3.545 1.12 3.485 1.12 3.485 1.44 3.365 1.44 3.365 1 3.425 1 3.425 0.5 2.22 0.5 2.22 0.6 1.695 0.6 1.695 1.46 1.575 1.46 1.575 0.6 1.095 0.6 1.095 1 1.155 1 1.155 1.24 0.975 1.24 0.975 0.9 0.24 0.9 0.24 1.64 0.355 1.64 0.355 1.88 0.235 1.88 0.235 1.76 0.12 1.76 0.12 0.78 0.135 0.78 0.135 0.66 0.255 0.66 0.255 0.78 0.975 0.78 0.975 0.48 2.1 0.48 2.1 0.38 3.765 0.38 3.765 0.36 4.005 0.36 ;
      POLYGON 3.005 1.22 2.855 1.22 2.855 1.62 2.915 1.62 2.915 1.74 2.675 1.74 2.675 1.62 2.735 1.62 2.735 1.16 2.075 1.16 2.075 1.18 1.835 1.18 1.835 1.04 2.735 1.04 2.735 0.72 2.975 0.72 2.975 0.84 2.855 0.84 2.855 0.98 3.005 0.98 ;
  END
END DFFSX2

MACRO DFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX2 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 1.31 0.935 1.55 ;
        RECT 0.595 1.52 0.855 1.67 ;
        RECT 0.735 1.43 0.935 1.55 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5 0.805 5.15 1.145 ;
        RECT 4.955 0.92 5.075 1.26 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.58 0.885 5.73 1.145 ;
        RECT 5.595 0.68 5.715 2.03 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.555 0.68 6.675 0.97 ;
        RECT 6.435 0.85 6.555 2.03 ;
        RECT 6.16 0.97 6.555 1.09 ;
        RECT 6.16 0.885 6.31 1.145 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.035 -0.18 7.155 0.73 ;
        RECT 6.015 -0.18 6.255 0.32 ;
        RECT 5.055 -0.18 5.295 0.32 ;
        RECT 3.735 -0.18 3.855 0.82 ;
        RECT 2.115 -0.18 2.355 0.32 ;
        RECT 0.675 -0.18 0.795 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.855 1.38 6.975 2.79 ;
        RECT 6.015 1.38 6.135 2.79 ;
        RECT 5.175 1.38 5.295 2.79 ;
        RECT 3.755 2.13 3.995 2.25 ;
        RECT 3.755 2.13 3.875 2.79 ;
        RECT 2.015 2.17 2.255 2.29 ;
        RECT 2.015 2.17 2.135 2.79 ;
        RECT 0.615 1.79 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.755 0.86 7.635 0.86 7.635 1.21 7.455 1.21 7.455 1.62 7.335 1.62 7.335 1.21 6.675 1.21 6.675 1.09 7.515 1.09 7.515 0.74 7.755 0.74 ;
      POLYGON 7.535 0.52 7.395 0.52 7.395 0.97 6.795 0.97 6.795 0.56 5.995 0.56 5.995 1.24 5.875 1.24 5.875 0.56 5.435 0.56 5.435 1.24 5.315 1.24 5.315 0.56 4.275 0.56 4.275 0.8 4.555 0.8 4.555 1.45 4.475 1.45 4.475 1.77 4.235 1.77 4.235 1.65 4.355 1.65 4.355 1.45 3.735 1.45 3.735 1.33 4.435 1.33 4.435 0.92 4.155 0.92 4.155 0.44 6.915 0.44 6.915 0.85 7.275 0.85 7.275 0.4 7.535 0.4 ;
      POLYGON 4.815 2.01 3.535 2.01 3.535 2.05 3.075 2.05 3.075 2.25 2.835 2.25 2.835 2.05 1.895 2.05 1.895 2.25 1.455 2.25 1.455 2.13 1.775 2.13 1.775 1.93 3.415 1.93 3.415 1.89 4.695 1.89 4.695 1.62 4.675 1.62 4.675 0.68 4.795 0.68 4.795 1.5 4.815 1.5 ;
      POLYGON 4.315 1.2 4.075 1.2 4.075 1.17 3.615 1.17 3.615 1.77 3.295 1.77 3.295 1.81 3.055 1.81 3.055 1.69 3.175 1.69 3.175 1.65 3.495 1.65 3.495 1.17 3.035 1.17 3.035 0.68 3.155 0.68 3.155 1.05 4.195 1.05 4.195 1.08 4.315 1.08 ;
      POLYGON 3.375 1.53 3.255 1.53 3.255 1.41 2.795 1.41 2.795 1.28 2.715 1.28 2.715 1.04 2.795 1.04 2.795 0.56 1.235 0.56 1.235 1.37 1.355 1.37 1.355 1.49 1.115 1.49 1.115 1.16 0.375 1.16 0.375 1.75 0.255 1.75 0.255 1.87 0.135 1.87 0.135 1.63 0.255 1.63 0.255 0.68 0.375 0.68 0.375 1.04 1.115 1.04 1.115 0.44 1.555 0.44 1.555 0.42 1.795 0.42 1.795 0.44 2.915 0.44 2.915 1.29 3.375 1.29 ;
      POLYGON 2.735 1.81 2.495 1.81 2.495 1.52 1.895 1.52 1.895 1.49 1.775 1.49 1.775 1.37 2.015 1.37 2.015 1.4 2.475 1.4 2.475 0.8 2.555 0.8 2.555 0.68 2.675 0.68 2.675 0.92 2.595 0.92 2.595 1.4 2.615 1.4 2.615 1.69 2.735 1.69 ;
      POLYGON 2.355 1.25 1.595 1.25 1.595 1.75 1.435 1.75 1.435 1.87 1.315 1.87 1.315 1.63 1.475 1.63 1.475 0.68 1.595 0.68 1.595 1.13 2.355 1.13 ;
  END
END DFFX2

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.795 0.24 1.22 ;
        RECT 0.07 0.795 0.24 1.2 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.625 0.675 1.99 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
        RECT 0.135 -0.18 0.255 0.675 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
END INVX1

MACRO OR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X6 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.67 0.82 2.79 1.17 ;
        RECT 0.39 0.82 2.79 0.94 ;
        RECT 0.39 0.82 0.51 1.15 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.06 2.39 1.3 ;
        RECT 2.1 1.06 2.25 1.435 ;
        RECT 1.03 1.06 2.39 1.18 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.3 1.79 1.42 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.55 1.3 1.67 1.725 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.49 0.93 5.35 1.05 ;
        RECT 5.23 0.4 5.35 1.05 ;
        RECT 5.03 1.41 5.15 2.21 ;
        RECT 3.35 1.41 5.15 1.53 ;
        RECT 4.41 0.885 4.57 1.145 ;
        RECT 4.41 0.795 4.53 1.53 ;
        RECT 4.39 0.4 4.51 1.05 ;
        RECT 4.19 1.41 4.31 2.21 ;
        RECT 3.49 0.4 3.61 1.05 ;
        RECT 3.35 1.41 3.47 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.81 -0.18 4.93 0.81 ;
        RECT 3.97 -0.18 4.09 0.81 ;
        RECT 2.95 0.34 3.19 0.46 ;
        RECT 2.95 -0.18 3.07 0.46 ;
        RECT 1.99 0.34 2.23 0.46 ;
        RECT 1.99 -0.18 2.11 0.46 ;
        RECT 1.03 0.34 1.27 0.46 ;
        RECT 1.03 -0.18 1.15 0.46 ;
        RECT 0.19 -0.18 0.31 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.61 1.65 4.73 2.79 ;
        RECT 3.77 1.65 3.89 2.79 ;
        RECT 2.93 1.795 3.05 2.79 ;
        RECT 0.61 1.56 0.73 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.29 1.29 3.03 1.29 3.03 1.675 1.91 1.675 1.91 2.21 1.79 2.21 1.79 1.555 2.91 1.555 2.91 0.7 0.55 0.7 0.55 0.58 3.03 0.58 3.03 1.17 4.29 1.17 ;
  END
END OR3X6

MACRO ADDFHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHXL 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.14 0.87 6.235 0.99 ;
        RECT 4.14 0.8 4.26 1.06 ;
        RECT 4.115 0.87 6.235 0.92 ;
        RECT 3.75 0.78 4.235 0.9 ;
        RECT 2.935 0.75 3.87 0.87 ;
        RECT 2.915 0.65 3.175 0.8 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.975 1.23 7.235 1.38 ;
        RECT 4.835 1.11 7.215 1.23 ;
        RECT 5.065 1.11 5.185 1.35 ;
        RECT 3.655 1.18 5.185 1.3 ;
        RECT 3.655 1.02 3.895 1.3 ;
        RECT 3.51 1.02 3.895 1.14 ;
        RECT 1.695 0.99 3.63 1.1 ;
        RECT 2.49 1.02 3.895 1.11 ;
        RECT 1.695 0.98 2.61 1.1 ;
        RECT 1.695 0.98 1.815 1.24 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.305 1.35 6.855 1.47 ;
        RECT 4.775 1.47 5.425 1.59 ;
        RECT 3.32 1.42 4.895 1.54 ;
        RECT 3.32 1.26 3.485 1.54 ;
        RECT 2.915 1.26 3.485 1.38 ;
        RECT 2.055 1.24 3.175 1.34 ;
        RECT 2.915 1.23 3.175 1.38 ;
        RECT 2.175 1.26 3.485 1.36 ;
        RECT 2.055 1.22 2.295 1.34 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2408 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 1.365 0.68 2.125 ;
        RECT 0.07 0.885 0.68 1.005 ;
        RECT 0.56 0.625 0.68 1.005 ;
        RECT 0.1 1.365 0.68 1.485 ;
        RECT 0.1 0.885 0.22 1.485 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2408 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.715 1.465 8.05 1.725 ;
        RECT 7.715 0.5 7.835 2.21 ;
    END
  END S
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.175 0.39 7.415 0.51 ;
        RECT 7.175 -0.18 7.295 0.51 ;
        RECT 4.835 0.39 5.075 0.51 ;
        RECT 4.835 -0.18 4.955 0.51 ;
        RECT 3.995 -0.18 4.115 0.64 ;
        RECT 1.715 -0.18 1.955 0.38 ;
        RECT 0.14 -0.18 0.26 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.175 2.07 7.415 2.19 ;
        RECT 7.175 2.07 7.295 2.79 ;
        RECT 4.825 2.29 5.065 2.79 ;
        RECT 3.865 1.9 3.985 2.79 ;
        RECT 3.745 1.9 3.985 2.15 ;
        RECT 1.715 2.22 1.955 2.79 ;
        RECT 0.14 1.605 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.595 1.55 7.475 1.55 7.475 1.95 6.295 1.95 6.295 2.21 6.175 2.21 6.175 1.95 5.905 1.95 5.905 2.17 5.785 2.17 5.785 1.83 7.355 1.83 7.355 0.75 5.795 0.75 5.795 0.49 5.915 0.49 5.915 0.63 6.315 0.63 6.315 0.49 6.435 0.49 6.435 0.63 7.475 0.63 7.475 1.43 7.595 1.43 ;
      POLYGON 6.085 1.71 5.665 1.71 5.665 2.17 4.105 2.17 4.105 1.78 3.55 1.78 3.55 2 3.285 2 3.285 2.21 3.165 2.21 3.165 2 2.795 2 2.795 2.1 0.995 2.1 0.995 1.245 0.34 1.245 0.34 1.125 0.995 1.125 0.995 0.5 2.675 0.5 2.675 0.41 3.415 0.41 3.415 0.46 3.535 0.46 3.535 0.58 3.295 0.58 3.295 0.53 2.795 0.53 2.795 0.82 2.675 0.82 2.675 0.62 1.115 0.62 1.115 1.98 2.675 1.98 2.675 1.48 2.795 1.48 2.795 1.88 3.165 1.88 3.165 1.69 3.285 1.69 3.285 1.88 3.43 1.88 3.43 1.66 4.225 1.66 4.225 2.05 5.545 2.05 5.545 1.59 6.085 1.59 ;
      POLYGON 5.495 0.75 4.475 0.75 4.475 0.68 4.355 0.68 4.355 0.56 4.595 0.56 4.595 0.63 5.375 0.63 5.375 0.5 5.495 0.5 ;
      POLYGON 5.425 1.89 5.185 1.89 5.185 1.86 4.585 1.86 4.585 1.93 4.345 1.93 4.345 1.74 5.185 1.74 5.185 1.71 5.425 1.71 ;
      RECT 1.235 0.74 2.435 0.86 ;
      POLYGON 2.375 1.86 2.255 1.86 2.255 1.6 1.535 1.6 1.535 1.86 1.415 1.86 1.415 1.34 1.535 1.34 1.535 1.48 2.375 1.48 ;
  END
END ADDFHXL

MACRO OAI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X2 0 0 ;
  SIZE 5.22 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.16 0.85 4.28 1.44 ;
        RECT 4.13 0.85 4.28 1.305 ;
    END
  END C0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.055 1.14 3.295 1.33 ;
        RECT 2.915 1.165 3.175 1.38 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.165 1.435 1.38 ;
        RECT 1.055 1.16 1.295 1.35 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.675 1.5 3.76 1.62 ;
        RECT 3.55 1.22 3.76 1.62 ;
        RECT 3.55 1.175 3.7 1.62 ;
        RECT 2.675 1.22 2.795 1.62 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.5 1.69 1.62 ;
        RECT 1.57 1.22 1.69 1.62 ;
        RECT 0.68 1.175 0.8 1.62 ;
        RECT 0.65 1.175 0.8 1.435 ;
        RECT 0.53 1.3 0.8 1.42 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7616 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.4 1.175 4.57 1.435 ;
        RECT 4.42 0.68 4.54 0.92 ;
        RECT 1.09 1.74 4.52 1.86 ;
        RECT 4.22 1.56 4.52 1.86 ;
        RECT 4.4 0.8 4.52 1.86 ;
        RECT 4.22 1.56 4.34 2.21 ;
        RECT 3.16 1.74 3.28 2.21 ;
        RECT 1.09 1.74 1.21 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.22 0.18 ;
        RECT 1.93 -0.18 2.05 0.73 ;
        RECT 1.09 -0.18 1.21 0.73 ;
        RECT 0.25 -0.18 0.37 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.22 2.79 ;
        RECT 4.64 1.56 4.76 2.79 ;
        RECT 3.74 1.98 3.98 2.15 ;
        RECT 3.74 1.98 3.86 2.79 ;
        RECT 1.67 1.98 1.91 2.15 ;
        RECT 1.67 1.98 1.79 2.79 ;
        RECT 0.45 1.74 0.57 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.96 0.73 4.84 0.73 4.84 0.56 4.12 0.56 4.12 0.73 4 0.73 4 0.56 3.28 0.56 3.28 0.73 3.16 0.73 3.16 0.56 2.44 0.56 2.44 0.73 2.32 0.73 2.32 0.44 4.96 0.44 ;
      POLYGON 3.76 0.86 3.64 0.86 3.64 0.97 0.67 0.97 0.67 0.68 0.79 0.68 0.79 0.85 1.51 0.85 1.51 0.68 1.63 0.68 1.63 0.85 2.74 0.85 2.74 0.68 2.86 0.68 2.86 0.85 3.52 0.85 3.52 0.74 3.76 0.74 ;
  END
END OAI221X2

MACRO SEDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX2 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.37 0.76 1.49 1.15 ;
        RECT 0.63 0.76 1.49 0.88 ;
        RECT 0.305 1.23 0.75 1.35 ;
        RECT 0.63 0.76 0.75 1.35 ;
        RECT 0.305 1.23 0.565 1.38 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.03 1.09 1.5 ;
        RECT 0.95 1 1.07 1.5 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.21 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 1.03 4.58 1.48 ;
        RECT 4.42 1.03 4.58 1.46 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.08 1.08 11.275 1.435 ;
        RECT 11.08 1.075 11.24 1.435 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.03 1.58 5.34 1.7 ;
        RECT 5 0.68 5.24 0.8 ;
        RECT 5.03 0.68 5.15 1.7 ;
        RECT 5 0.68 5.15 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.76 -0.18 10.88 0.715 ;
        RECT 8.77 -0.18 9.01 0.39 ;
        RECT 6.97 0.46 7.21 0.58 ;
        RECT 6.97 -0.18 7.09 0.58 ;
        RECT 5.48 -0.18 5.72 0.32 ;
        RECT 4.52 -0.18 4.64 0.67 ;
        RECT 2.35 0.46 2.59 0.58 ;
        RECT 2.35 -0.18 2.47 0.58 ;
        RECT 0.87 -0.18 0.99 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 10.8 1.795 10.92 2.79 ;
        RECT 8.57 2.25 8.81 2.79 ;
        RECT 6.85 1.47 6.97 2.79 ;
        RECT 5.58 2.06 5.82 2.18 ;
        RECT 5.58 2.06 5.7 2.79 ;
        RECT 4.74 2.06 4.86 2.79 ;
        RECT 4.62 2.06 4.86 2.18 ;
        RECT 2.41 1.57 2.53 2.79 ;
        RECT 0.81 1.86 0.93 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.4 1.855 11.16 1.855 11.16 1.675 10.68 1.675 10.68 2.25 9.13 2.25 9.13 2.13 8.19 2.13 8.19 2.25 7.83 2.25 7.83 2.13 8.07 2.13 8.07 2.01 9.355 2.01 9.355 2.13 10.56 2.13 10.56 1.555 10.84 1.555 10.84 0.955 10.72 0.955 10.72 1.075 10.6 1.075 10.6 0.835 11.18 0.835 11.18 0.475 11.3 0.475 11.3 0.955 10.96 0.955 10.96 1.555 11.28 1.555 11.28 1.735 11.4 1.735 ;
      POLYGON 10.46 0.715 10.44 0.715 10.44 2.01 9.63 2.01 9.63 1.89 7.85 1.89 7.85 1.33 7.45 1.33 7.45 1.21 7.85 1.21 7.85 0.99 8.27 0.99 8.27 1.11 7.97 1.11 7.97 1.77 9.63 1.77 9.63 1.33 9.53 1.33 9.53 1.21 9.77 1.21 9.77 1.33 9.75 1.33 9.75 1.89 10.32 1.89 10.32 0.595 10.34 0.595 10.34 0.475 10.46 0.475 ;
      POLYGON 10.11 1.77 9.87 1.77 9.87 1.53 9.95 1.53 9.95 0.48 9.25 0.48 9.25 0.63 8.53 0.63 8.53 0.48 7.49 0.48 7.49 0.82 6.73 0.82 6.73 0.53 6.055 0.53 6.055 0.56 4.88 0.56 4.88 0.91 4.145 0.91 4.145 0.86 4 0.86 4 1.77 3.88 1.77 3.88 0.62 4 0.62 4 0.74 4.265 0.74 4.265 0.79 4.76 0.79 4.76 0.44 5.935 0.44 5.935 0.41 6.85 0.41 6.85 0.7 7.37 0.7 7.37 0.36 8.65 0.36 8.65 0.51 9.13 0.51 9.13 0.36 10.07 0.36 10.07 1.53 10.11 1.53 ;
      POLYGON 9.71 0.72 9.59 0.72 9.59 1.09 9.41 1.09 9.41 1.53 9.51 1.53 9.51 1.65 9.27 1.65 9.27 1.53 9.29 1.53 9.29 1.36 8.63 1.36 8.63 1.12 8.75 1.12 8.75 1.24 9.29 1.24 9.29 0.97 9.47 0.97 9.47 0.6 9.71 0.6 ;
      POLYGON 9.07 1.12 8.95 1.12 8.95 1 8.51 1 8.51 1.65 8.09 1.65 8.09 1.53 8.39 1.53 8.39 0.87 8.17 0.87 8.17 0.6 8.41 0.6 8.41 0.75 8.51 0.75 8.51 0.88 9.07 0.88 ;
      POLYGON 7.99 0.72 7.73 0.72 7.73 1.06 7.33 1.06 7.33 1.45 7.73 1.45 7.73 1.99 7.61 1.99 7.61 1.57 7.21 1.57 7.21 1.35 6.61 1.35 6.61 1.33 6.49 1.33 6.49 1.21 6.73 1.21 6.73 1.23 7.21 1.23 7.21 0.94 7.61 0.94 7.61 0.6 7.99 0.6 ;
      POLYGON 7.09 1.11 6.85 1.11 6.85 1.09 6.37 1.09 6.37 1.47 6.55 1.47 6.55 1.78 6.43 1.78 6.43 1.59 6.25 1.59 6.25 1.21 6.18 1.21 6.18 0.97 6.25 0.97 6.25 0.92 6.37 0.92 6.37 0.65 6.61 0.65 6.61 0.97 6.97 0.97 6.97 0.99 7.09 0.99 ;
      POLYGON 6.24 2.17 6.12 2.17 6.12 2.05 5.94 2.05 5.94 1.94 4.48 1.94 4.48 2.25 2.65 2.25 2.65 1.45 2.27 1.45 2.27 1.21 2.39 1.21 2.39 1.33 2.77 1.33 2.77 2.13 4.36 2.13 4.36 1.82 5.94 1.82 5.94 0.68 6.2 0.68 6.2 0.8 6.06 0.8 6.06 1.82 6.24 1.82 ;
      POLYGON 4.24 2.01 2.89 2.01 2.89 1.33 3.005 1.33 3.005 0.77 2.95 0.77 2.95 0.65 3.19 0.65 3.19 0.77 3.125 0.77 3.125 1.45 3.01 1.45 3.01 1.89 3.64 1.89 3.64 1.2 3.56 1.2 3.56 0.96 3.76 0.96 3.76 1.89 4.12 1.89 4.12 1.2 4.24 1.2 ;
      POLYGON 3.52 0.77 3.44 0.77 3.44 1.52 3.52 1.52 3.52 1.77 3.4 1.77 3.4 1.64 3.32 1.64 3.32 0.65 3.4 0.65 3.4 0.53 2.83 0.53 2.83 0.82 1.77 0.82 1.77 0.83 1.73 0.83 1.73 1.66 1.57 1.66 1.57 2.01 1.45 2.01 1.45 1.54 1.61 1.54 1.61 0.71 1.65 0.71 1.65 0.59 1.77 0.59 1.77 0.7 2.71 0.7 2.71 0.41 3.52 0.41 ;
      POLYGON 2.09 1.09 1.97 1.09 1.97 2.25 1.21 2.25 1.21 1.74 0.45 1.74 0.45 1.86 0.33 1.86 0.33 1.74 0.065 1.74 0.065 0.99 0.39 0.99 0.39 0.59 0.51 0.59 0.51 1.11 0.185 1.11 0.185 1.62 1.21 1.62 1.21 1.3 1.49 1.3 1.49 1.42 1.33 1.42 1.33 2.13 1.85 2.13 1.85 0.97 2.09 0.97 ;
  END
END SEDFFHQX2

MACRO SDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX1 0 0 ;
  SIZE 10.44 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.005 1.22 2.125 1.46 ;
        RECT 1.755 1.52 2.015 1.67 ;
        RECT 1.895 1.34 2.015 1.67 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.74 1.185 7.015 1.435 ;
        RECT 6.74 1.165 6.89 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.715 0.94 8.975 1.09 ;
        RECT 8.715 0.94 8.955 1.3 ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.165 9.555 1.38 ;
        RECT 9.215 0.98 9.335 1.36 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.775 0.885 10.08 1.22 ;
        RECT 9.93 0.88 10.08 1.22 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.99 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 2.21 ;
        RECT 1.23 0.885 1.485 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.44 0.18 ;
        RECT 9.075 -0.18 9.195 0.82 ;
        RECT 6.995 -0.18 7.115 0.84 ;
        RECT 4.885 -0.18 5.125 0.32 ;
        RECT 3.105 -0.18 3.345 0.32 ;
        RECT 1.785 -0.18 1.905 0.73 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.44 2.79 ;
        RECT 9.915 1.58 10.035 2.79 ;
        RECT 9.015 2.06 9.135 2.79 ;
        RECT 6.995 1.88 7.115 2.79 ;
        RECT 4.945 2.14 5.065 2.79 ;
        RECT 3.285 2.08 3.525 2.2 ;
        RECT 3.285 2.08 3.405 2.79 ;
        RECT 1.785 1.79 1.905 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.32 1.46 9.795 1.46 9.795 1.62 9.615 1.62 9.615 1.86 9.235 1.86 9.235 1.94 8.175 1.94 8.175 2 8.055 2 8.055 1.44 8.235 1.44 8.235 0.84 8.115 0.84 8.115 0.6 8.235 0.6 8.235 0.72 8.355 0.72 8.355 1.56 8.175 1.56 8.175 1.82 9.115 1.82 9.115 1.74 9.495 1.74 9.495 1.5 9.675 1.5 9.675 1.34 10.2 1.34 10.2 0.76 9.655 0.76 9.655 0.64 10.32 0.64 ;
      POLYGON 8.775 0.82 8.595 0.82 8.595 1.42 8.655 1.42 8.655 1.7 8.535 1.7 8.535 1.54 8.475 1.54 8.475 0.7 8.655 0.7 8.655 0.48 7.995 0.48 7.995 0.98 8.115 0.98 8.115 1.1 7.995 1.1 7.995 1.32 7.495 1.32 7.495 1.44 7.375 1.44 7.375 1.2 7.875 1.2 7.875 0.36 8.775 0.36 ;
      POLYGON 7.755 1.08 7.255 1.08 7.255 1.56 7.755 1.56 7.755 2 7.635 2 7.635 1.68 6.365 1.68 6.365 1.72 6.125 1.72 6.125 1.6 6.245 1.6 6.245 0.92 6.185 0.92 6.185 0.68 6.305 0.68 6.305 0.8 6.365 0.8 6.365 1.56 7.135 1.56 7.135 0.96 7.635 0.96 7.635 0.6 7.755 0.6 ;
      POLYGON 6.755 1.96 5.885 1.96 5.885 0.98 5.945 0.98 5.945 0.56 4.345 0.56 4.345 1.24 4.225 1.24 4.225 0.44 5.425 0.44 5.425 0.4 5.665 0.4 5.665 0.44 6.545 0.44 6.545 0.48 6.695 0.48 6.695 0.84 6.575 0.84 6.575 0.6 6.425 0.6 6.425 0.56 6.065 0.56 6.065 1.1 6.005 1.1 6.005 1.28 6.125 1.28 6.125 1.4 6.005 1.4 6.005 1.84 6.755 1.84 ;
      POLYGON 5.825 0.86 5.765 0.86 5.765 1.78 5.645 1.78 5.645 1.44 4.825 1.44 4.825 1.4 4.705 1.4 4.705 1.28 4.945 1.28 4.945 1.32 5.645 1.32 5.645 0.86 5.585 0.86 5.585 0.74 5.825 0.74 ;
      POLYGON 5.685 2.16 5.445 2.16 5.445 2.02 4.365 2.02 4.365 2.16 4.125 2.16 4.125 2.02 3.645 2.02 3.645 1.96 2.53 1.96 2.53 1.92 2.265 1.92 2.265 0.68 2.385 0.68 2.385 1.8 2.65 1.8 2.65 1.84 3.645 1.84 3.645 1.18 3.625 1.18 3.625 1.06 3.865 1.06 3.865 1.18 3.765 1.18 3.765 1.9 5.565 1.9 5.565 2.04 5.685 2.04 ;
      POLYGON 5.345 1.2 5.105 1.2 5.105 1.16 4.585 1.16 4.585 1.78 4.465 1.78 4.465 0.68 4.585 0.68 4.585 1.04 5.225 1.04 5.225 1.08 5.345 1.08 ;
      POLYGON 4.165 1.78 4.045 1.78 4.045 1.48 3.985 1.48 3.985 0.92 3.825 0.92 3.825 0.68 2.895 0.68 2.895 0.56 2.745 0.56 2.745 0.4 2.985 0.4 2.985 0.44 3.015 0.44 3.015 0.56 3.945 0.56 3.945 0.8 4.105 0.8 4.105 1.36 4.165 1.36 ;
      POLYGON 3.505 1.18 2.925 1.18 2.925 1.6 3.045 1.6 3.045 1.72 2.805 1.72 2.805 0.92 2.655 0.92 2.655 0.8 2.505 0.8 2.505 0.56 2.145 0.56 2.145 0.97 1.765 0.97 1.765 1.24 1.645 1.24 1.645 0.85 2.025 0.85 2.025 0.44 2.625 0.44 2.625 0.68 2.775 0.68 2.775 0.8 2.925 0.8 2.925 1.06 3.505 1.06 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END SDFFTRX1

MACRO AND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X2 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.225 0.565 1.495 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.09 1.44 ;
        RECT 0.805 1.175 1.09 1.345 ;
        RECT 0.805 1.1 0.925 1.345 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.225 1.015 1.38 1.47 ;
        RECT 1.225 1.015 1.345 1.495 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.105 1.96 1.435 ;
        RECT 1.74 1.09 1.86 1.415 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.32 0.885 2.54 1.145 ;
        RECT 2.32 0.61 2.44 1.48 ;
        RECT 2.225 1.36 2.345 2.08 ;
        RECT 2.22 0.49 2.34 0.73 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 2.64 -0.18 2.76 0.73 ;
        RECT 1.8 -0.18 1.92 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.645 1.43 2.765 2.79 ;
        RECT 1.805 1.555 1.925 2.79 ;
        RECT 1.025 2.195 1.145 2.79 ;
        RECT 0.135 2.195 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.2 1.24 2.08 1.24 2.08 0.97 1.62 0.97 1.62 1.735 1.505 1.735 1.505 1.855 1.385 1.855 1.385 1.735 0.485 1.735 0.485 1.615 1.5 1.615 1.5 0.86 0.265 0.86 0.265 0.74 1.62 0.74 1.62 0.85 2.2 0.85 ;
  END
END AND4X2

MACRO OAI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.36 1.38 1.725 ;
        RECT 1.21 1.28 1.33 1.65 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.165 1.67 1.62 ;
        RECT 1.53 1.1 1.65 1.62 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.08 0.51 1.53 ;
        RECT 0.36 1.08 0.48 1.555 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.98 0.82 1.405 ;
        RECT 0.65 1.175 0.8 1.585 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.28 0.86 1.58 0.98 ;
        RECT 1.46 0.68 1.58 0.98 ;
        RECT 0.97 1.04 1.4 1.16 ;
        RECT 1.28 0.86 1.4 1.16 ;
        RECT 0.97 1.04 1.09 1.86 ;
        RECT 0.94 1.465 1.09 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.69 1.74 1.81 2.79 ;
        RECT 0.22 1.74 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2 0.92 1.88 0.92 1.88 0.56 1.16 0.56 1.16 0.92 1.04 0.92 1.04 0.86 0.075 0.86 0.075 0.74 1.04 0.74 1.04 0.44 2 0.44 ;
  END
END OAI22XL

MACRO DFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX4 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 0.63 1.67 2.21 ;
        RECT 0.65 1.315 1.67 1.435 ;
        RECT 0.71 0.63 0.83 2.21 ;
        RECT 0.65 1.175 0.83 1.435 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.485 0.7 5.605 1.08 ;
        RECT 4.955 0.7 5.605 0.82 ;
        RECT 4.955 0.36 5.075 0.82 ;
        RECT 3.895 0.36 5.075 0.48 ;
        RECT 3.55 0.44 4.015 0.56 ;
        RECT 3.55 0.885 3.7 1.145 ;
        RECT 2.91 1.22 3.67 1.34 ;
        RECT 3.55 0.44 3.67 1.34 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.845 1.18 8.105 1.41 ;
        RECT 7.905 1.02 8.025 1.43 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.215 1.02 9.335 1.26 ;
        RECT 9.005 1.23 9.265 1.38 ;
        RECT 9.145 1.14 9.335 1.26 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.455 -0.18 9.575 0.92 ;
        RECT 7.925 0.54 8.165 0.66 ;
        RECT 7.925 -0.18 8.045 0.66 ;
        RECT 6.405 -0.18 6.525 0.69 ;
        RECT 5.265 0.46 5.505 0.58 ;
        RECT 5.385 -0.18 5.505 0.58 ;
        RECT 2.81 -0.18 2.93 0.68 ;
        RECT 1.97 -0.18 2.09 0.68 ;
        RECT 1.13 -0.18 1.25 0.68 ;
        RECT 0.29 -0.18 0.41 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.395 1.46 9.515 2.79 ;
        RECT 8.065 1.79 8.185 2.79 ;
        RECT 6.31 2.29 6.55 2.79 ;
        RECT 5.35 2.29 5.59 2.79 ;
        RECT 3.65 1.94 3.77 2.79 ;
        RECT 2.81 1.7 2.93 2.79 ;
        RECT 1.97 1.69 2.09 2.79 ;
        RECT 1.13 1.56 1.25 2.79 ;
        RECT 0.29 1.56 0.41 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.155 1.62 8.765 1.62 8.765 0.84 8.975 0.84 8.975 0.48 8.405 0.48 8.405 1.06 8.165 1.06 8.165 0.9 7.665 0.9 7.665 1.05 7.445 1.05 7.445 1.93 5.205 1.93 5.205 1.86 4.86 1.86 4.86 1.3 4.18 1.3 4.18 1.04 4.06 1.04 4.06 0.92 4.3 0.92 4.3 1.18 5.1 1.18 5.1 1.3 4.98 1.3 4.98 1.74 5.325 1.74 5.325 1.81 7.325 1.81 7.325 1.29 6.845 1.29 6.845 1.17 7.325 1.17 7.325 0.78 8.285 0.78 8.285 0.36 9.095 0.36 9.095 0.96 8.885 0.96 8.885 1.5 9.155 1.5 ;
      POLYGON 8.765 0.72 8.645 0.72 8.645 1.3 8.605 1.3 8.605 1.91 8.485 1.91 8.485 1.67 7.685 1.67 7.685 2.17 5.17 2.17 5.17 2.24 4.4 2.24 4.4 2.12 5.05 2.12 5.05 2.05 7.565 2.05 7.565 1.19 7.685 1.19 7.685 1.55 8.485 1.55 8.485 1.18 8.525 1.18 8.525 0.6 8.765 0.6 ;
      POLYGON 7.525 0.66 7.205 0.66 7.205 1.05 6.725 1.05 6.725 1.45 7.085 1.45 7.085 1.57 7.205 1.57 7.205 1.69 6.965 1.69 6.965 1.57 6.605 1.57 6.605 1.29 6.085 1.29 6.085 1.33 5.965 1.33 5.965 1.09 6.085 1.09 6.085 1.17 6.605 1.17 6.605 0.93 7.085 0.93 7.085 0.54 7.525 0.54 ;
      POLYGON 6.485 1.05 6.205 1.05 6.205 0.97 5.845 0.97 5.845 1.57 6.07 1.57 6.07 1.69 5.725 1.69 5.725 1.32 5.34 1.32 5.34 1.62 5.1 1.62 5.1 1.5 5.22 1.5 5.22 1.06 4.715 1.06 4.715 0.72 4.56 0.72 4.56 0.6 4.835 0.6 4.835 0.94 5.34 0.94 5.34 1.2 5.725 1.2 5.725 0.85 5.965 0.85 5.965 0.5 6.085 0.5 6.085 0.85 6.325 0.85 6.325 0.93 6.485 0.93 ;
      POLYGON 4.74 1.96 4.62 1.96 4.62 1.58 2.63 1.58 2.63 1.33 2.75 1.33 2.75 1.46 3.82 1.46 3.82 0.68 4.14 0.68 4.14 0.6 4.38 0.6 4.38 0.72 4.26 0.72 4.26 0.8 3.94 0.8 3.94 1.46 4.62 1.46 4.62 1.44 4.74 1.44 ;
      POLYGON 4.38 1.9 4.14 1.9 4.14 1.82 3.35 1.82 3.35 2.21 3.23 2.21 3.23 1.7 4.38 1.7 ;
      POLYGON 3.43 1.1 3.31 1.1 3.31 1.07 2.51 1.07 2.51 2.21 2.39 2.21 2.39 1.07 1.95 1.07 1.95 1.19 1.83 1.19 1.83 0.95 2.39 0.95 2.39 0.54 2.51 0.54 2.51 0.95 3.31 0.95 3.31 0.86 3.43 0.86 ;
  END
END DFFSHQX4

MACRO NOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2XL 0 0 ;
  SIZE 1.16 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.025 0.675 1.265 ;
        RECT 0.39 1.145 0.675 1.265 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.79 0.24 1.225 ;
        RECT 0.07 0.73 0.22 1.145 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.795 0.785 0.915 1.825 ;
        RECT 0.65 1.465 0.915 1.725 ;
        RECT 0.495 0.785 0.915 0.905 ;
        RECT 0.495 0.665 0.615 0.905 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.16 0.18 ;
        RECT 0.905 -0.18 1.025 0.385 ;
        RECT 0.135 -0.18 0.255 0.385 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.16 2.79 ;
        RECT 0.155 1.705 0.275 2.79 ;
    END
  END VDD
END NOR2XL

MACRO XNOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X2 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.11 1.725 1.38 ;
        RECT 1.465 1.02 1.705 1.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.26 3.525 1.38 ;
        RECT 2.625 1.23 2.885 1.38 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 1.175 1.09 1.435 ;
        RECT 0.665 1.62 0.945 1.74 ;
        RECT 0.825 0.68 0.945 1.74 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.125 0.72 3.365 0.84 ;
        RECT 3.205 -0.18 3.325 0.84 ;
        RECT 1.245 -0.18 1.365 0.73 ;
        RECT 0.405 -0.18 0.525 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 3.125 1.74 3.365 1.86 ;
        RECT 3.125 1.74 3.245 2.79 ;
        RECT 1.145 2.1 1.385 2.22 ;
        RECT 1.145 2.1 1.265 2.79 ;
        RECT 0.185 2.1 0.425 2.22 ;
        RECT 0.185 2.1 0.305 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.765 1.68 3.725 1.68 3.725 1.8 3.605 1.8 3.605 1.62 2.655 1.62 2.655 2.22 1.885 2.22 1.885 2.1 2.535 2.1 2.535 1.5 3.645 1.5 3.645 1.11 2.505 1.11 2.505 1.24 2.385 1.24 2.385 0.99 3.605 0.99 3.605 0.66 3.725 0.66 3.725 0.87 3.765 0.87 ;
      POLYGON 3.085 0.52 1.905 0.52 1.905 0.66 1.845 0.66 1.845 0.78 1.965 0.78 1.965 1.74 1.625 1.74 1.625 1.62 1.845 1.62 1.845 0.9 1.725 0.9 1.725 0.54 1.785 0.54 1.785 0.4 3.085 0.4 ;
      POLYGON 2.265 1.98 0.425 1.98 0.425 1.36 0.545 1.36 0.545 1.24 0.665 1.24 0.665 1.48 0.545 1.48 0.545 1.86 2.145 1.86 2.145 0.66 2.265 0.66 ;
  END
END XNOR2X2

MACRO SEDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX2 0 0 ;
  SIZE 12.76 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.905 1.28 7.025 1.52 ;
        RECT 6.74 1.28 7.025 1.435 ;
        RECT 6.74 1.175 6.89 1.435 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.23 7.525 1.445 ;
        RECT 7.325 1.23 7.445 1.64 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.18 9.555 1.45 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.615 1.21 11.915 1.425 ;
        RECT 11.615 1.21 11.875 1.45 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 1.23 12.455 1.38 ;
        RECT 12.165 1.21 12.315 1.33 ;
        RECT 12.165 0.97 12.285 1.33 ;
        RECT 11.045 0.97 12.285 1.09 ;
        RECT 11.045 0.97 11.495 1.17 ;
        RECT 11.045 0.97 11.165 1.77 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 0.68 0.675 1.99 ;
        RECT 0.36 0.885 0.675 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.945 1.465 10.185 1.74 ;
        RECT 10.065 0.67 10.185 1.74 ;
        RECT 9.93 1.465 10.185 1.725 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.76 0.18 ;
        RECT 11.815 0.73 12.055 0.85 ;
        RECT 11.815 -0.18 11.935 0.85 ;
        RECT 10.545 -0.18 10.665 0.39 ;
        RECT 9.585 0.54 9.825 0.66 ;
        RECT 9.705 -0.18 9.825 0.66 ;
        RECT 7.165 -0.18 7.285 0.8 ;
        RECT 5.54 -0.18 5.66 0.9 ;
        RECT 3.4 0.61 3.64 0.73 ;
        RECT 3.52 -0.18 3.64 0.73 ;
        RECT 1.8 -0.18 1.92 0.53 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.76 2.79 ;
        RECT 11.905 1.97 12.025 2.79 ;
        RECT 10.425 2.1 10.665 2.22 ;
        RECT 10.425 2.1 10.545 2.79 ;
        RECT 9.465 2.1 9.705 2.22 ;
        RECT 9.465 2.1 9.585 2.79 ;
        RECT 7.265 2.24 7.505 2.79 ;
        RECT 5.54 1.88 5.66 2.79 ;
        RECT 5.42 1.88 5.66 2 ;
        RECT 3.52 1.81 3.64 2.79 ;
        RECT 3.4 1.81 3.64 1.93 ;
        RECT 1.64 2.01 1.76 2.79 ;
        RECT 1.035 2.14 1.155 2.79 ;
        RECT 0.135 1.34 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.695 1.97 12.445 1.97 12.445 2.09 12.325 2.09 12.325 1.85 12.575 1.85 12.575 1.69 11.345 1.69 11.345 1.57 12.575 1.57 12.575 0.85 12.235 0.85 12.235 0.73 12.695 0.73 ;
      POLYGON 11.415 0.85 10.925 0.85 10.925 1.91 11.365 1.91 11.365 2.03 10.805 2.03 10.805 1.98 8.445 1.98 8.445 1.62 8.745 1.62 8.745 0.74 8.165 0.74 8.165 0.62 8.865 0.62 8.865 1.74 8.565 1.74 8.565 1.86 10.805 1.86 10.805 0.73 11.415 0.73 ;
      POLYGON 9.905 1.23 9.785 1.23 9.785 0.9 9.345 0.9 9.345 0.5 7.525 0.5 7.525 1.04 6.925 1.04 6.925 0.5 6.25 0.5 6.25 0.66 6.08 0.66 6.08 0.9 6.38 0.9 6.38 1.58 6.26 1.58 6.26 1.02 5.96 1.02 5.96 0.54 6.13 0.54 6.13 0.38 7.045 0.38 7.045 0.92 7.405 0.92 7.405 0.38 9.465 0.38 9.465 0.78 9.905 0.78 ;
      POLYGON 9.225 0.74 9.105 0.74 9.105 0.94 9.225 0.94 9.225 1.06 9.105 1.06 9.105 1.62 9.225 1.62 9.225 1.74 8.985 1.74 8.985 0.62 9.225 0.62 ;
      POLYGON 8.625 1.5 7.885 1.5 7.885 1.38 8.505 1.38 8.505 0.9 8.625 0.9 ;
      POLYGON 8.145 1.88 8.025 1.88 8.025 1.76 7.765 1.76 7.765 1.88 7.235 1.88 7.235 2.12 6.32 2.12 6.32 2.06 5.78 2.06 5.78 1.76 4.84 1.76 4.84 1.77 4.7 1.77 4.7 1.89 4.58 1.89 4.58 1.65 4.7 1.65 4.7 0.62 4.82 0.62 4.82 1.64 5.9 1.64 5.9 1.94 6.44 1.94 6.44 2 7.115 2 7.115 1.76 7.645 1.76 7.645 1.14 7.745 1.14 7.745 0.62 7.985 0.62 7.985 0.74 7.865 0.74 7.865 1.26 7.765 1.26 7.765 1.64 8.145 1.64 ;
      POLYGON 6.965 1.88 6.845 1.88 6.845 1.82 6.02 1.82 6.02 1.52 5.81 1.52 5.81 1.26 5.28 1.26 5.28 1.02 5.4 1.02 5.4 1.14 5.93 1.14 5.93 1.4 6.14 1.4 6.14 1.7 6.5 1.7 6.5 0.62 6.805 0.62 6.805 0.74 6.62 0.74 6.62 1.64 6.965 1.64 ;
      POLYGON 5.3 2.2 3.76 2.2 3.76 1.69 3.28 1.69 3.28 2.11 2.16 2.11 2.16 2.25 1.92 2.25 1.92 2.13 2.04 2.13 2.04 1.89 1.66 1.89 1.66 1.84 1.395 1.84 1.395 1.46 1.215 1.46 1.215 1.2 0.795 1.2 0.795 1.08 1.215 1.08 1.215 0.74 1.635 0.74 1.635 0.86 1.335 0.86 1.335 1.34 1.515 1.34 1.515 1.72 1.78 1.72 1.78 1.77 2.16 1.77 2.16 1.99 3.16 1.99 3.16 1.57 3.88 1.57 3.88 2.08 5.3 2.08 ;
      POLYGON 5.24 0.9 5.16 0.9 5.16 1.4 5.18 1.4 5.18 1.52 4.94 1.52 4.94 1.4 5.04 1.4 5.04 0.78 5.12 0.78 5.12 0.66 4.94 0.66 4.94 0.5 4.58 0.5 4.58 1.04 4.56 1.04 4.56 1.53 4.44 1.53 4.44 0.92 4.46 0.92 4.46 0.5 3.88 0.5 3.88 0.97 3.16 0.97 3.16 0.5 2.32 0.5 2.32 1.29 2.4 1.29 2.4 1.41 2.16 1.41 2.16 1.29 2.2 1.29 2.2 0.38 2.61 0.38 2.61 0.36 2.85 0.36 2.85 0.38 3.28 0.38 3.28 0.85 3.76 0.85 3.76 0.38 3.96 0.38 3.96 0.36 4.2 0.36 4.2 0.38 5.06 0.38 5.06 0.54 5.24 0.54 ;
      POLYGON 4.34 0.8 4.22 0.8 4.22 1.63 4.28 1.63 4.28 1.87 4.16 1.87 4.16 1.75 4.1 1.75 4.1 1.21 3.18 1.21 3.18 1.09 4.1 1.09 4.1 0.68 4.34 0.68 ;
      POLYGON 3.84 1.45 3.04 1.45 3.04 1.87 2.92 1.87 2.92 0.62 3.04 0.62 3.04 1.33 3.84 1.33 ;
      POLYGON 2.68 0.8 2.64 0.8 2.64 1.69 2.68 1.69 2.68 1.81 2.44 1.81 2.44 1.65 1.9 1.65 1.9 1.2 1.455 1.2 1.455 1.08 2.02 1.08 2.02 1.53 2.52 1.53 2.52 0.8 2.44 0.8 2.44 0.68 2.68 0.68 ;
  END
END SEDFFX2

MACRO NAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X8 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.855 1.05 5.095 1.17 ;
        RECT 0.305 0.965 4.975 1.085 ;
        RECT 3.695 0.965 3.935 1.17 ;
        RECT 1.815 0.965 2.055 1.17 ;
        RECT 0.435 0.965 0.675 1.175 ;
        RECT 0.305 0.94 0.565 1.09 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.375 1.19 5.835 1.31 ;
        RECT 1.175 1.29 5.495 1.41 ;
        RECT 5.235 1.23 5.835 1.31 ;
        RECT 4.055 1.21 4.295 1.41 ;
        RECT 2.875 1.205 3.115 1.41 ;
        RECT 1.055 1.205 1.295 1.325 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.2732 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.53 6.075 1.65 ;
        RECT 5.955 0.71 6.075 1.65 ;
        RECT 5.87 1.465 6.02 1.725 ;
        RECT 0.915 0.71 6.075 0.83 ;
        RECT 5.595 1.53 5.715 2.21 ;
        RECT 4.755 1.53 4.875 2.21 ;
        RECT 3.915 1.53 4.035 2.21 ;
        RECT 3.075 1.53 3.195 2.21 ;
        RECT 2.235 1.53 2.355 2.21 ;
        RECT 1.395 1.53 1.515 2.21 ;
        RECT 0.555 1.465 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.115 0.46 5.355 0.58 ;
        RECT 5.115 -0.18 5.235 0.58 ;
        RECT 3.555 0.46 3.795 0.58 ;
        RECT 3.555 -0.18 3.675 0.58 ;
        RECT 1.555 0.46 1.795 0.58 ;
        RECT 1.555 -0.18 1.675 0.58 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 6.015 1.845 6.135 2.79 ;
        RECT 5.175 1.77 5.295 2.79 ;
        RECT 4.335 1.77 4.455 2.79 ;
        RECT 3.495 1.77 3.615 2.79 ;
        RECT 2.655 1.77 2.775 2.79 ;
        RECT 1.815 1.77 1.935 2.79 ;
        RECT 0.975 1.77 1.095 2.79 ;
        RECT 0.135 1.465 0.255 2.79 ;
    END
  END VDD
END NAND2X8

MACRO SDFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX4 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.915 0.72 2.155 0.84 ;
        RECT 1.935 1.28 2.055 2.04 ;
        RECT 1.915 0.72 2.035 1.4 ;
        RECT 0.94 1.025 2.035 1.145 ;
        RECT 1.095 0.72 1.215 2.04 ;
        RECT 0.94 0.885 1.215 1.145 ;
        RECT 0.955 0.72 1.215 1.145 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.475 0.98 0.8 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
        RECT 0.475 0.98 0.595 1.22 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.16 7.525 1.38 ;
        RECT 7.385 1.12 7.505 1.51 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 1.22 8.745 1.44 ;
        RECT 8.425 1.22 8.685 1.465 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.885 0.98 9.065 1.1 ;
        RECT 8.715 0.94 8.975 1.1 ;
        RECT 7.645 1.39 8.005 1.51 ;
        RECT 7.885 0.98 8.005 1.51 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.725 -0.18 8.845 0.82 ;
        RECT 7.265 0.64 7.505 0.76 ;
        RECT 7.385 -0.18 7.505 0.76 ;
        RECT 5.175 -0.18 5.295 0.38 ;
        RECT 3.475 -0.18 3.595 0.38 ;
        RECT 2.395 -0.18 2.635 0.36 ;
        RECT 1.435 -0.18 1.675 0.36 ;
        RECT 0.475 -0.18 0.595 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.565 1.93 8.805 2.05 ;
        RECT 8.565 1.93 8.685 2.79 ;
        RECT 7.225 1.87 7.345 2.79 ;
        RECT 4.935 2.2 5.175 2.79 ;
        RECT 3.255 1.66 3.375 2.79 ;
        RECT 2.355 1.39 2.475 2.79 ;
        RECT 1.515 1.39 1.635 2.79 ;
        RECT 0.675 1.39 0.795 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.305 1.825 9.165 1.825 9.165 1.99 9.045 1.99 9.045 1.705 8.125 1.705 8.125 1.43 8.245 1.43 8.245 1.585 9.185 1.585 9.185 0.82 9.145 0.82 9.145 0.58 9.265 0.58 9.265 0.7 9.305 0.7 ;
      POLYGON 8.205 0.82 7.765 0.82 7.765 1 7.145 1 7.145 1.63 7.985 1.63 7.985 1.99 7.865 1.99 7.865 1.75 6.375 1.75 6.375 1.9 6.255 1.9 6.255 1.63 7.025 1.63 7.025 0.52 6.515 0.52 6.515 0.84 6.275 0.84 6.275 0.72 6.395 0.72 6.395 0.4 7.145 0.4 7.145 0.88 7.645 0.88 7.645 0.7 8.085 0.7 8.085 0.58 8.205 0.58 ;
      POLYGON 6.985 2.05 6.865 2.05 6.865 2.14 6.015 2.14 6.015 2.08 4.215 2.08 4.215 1.44 4.035 1.44 4.035 1.56 3.915 1.56 3.915 1.32 4.215 1.32 4.215 1.12 4.455 1.12 4.455 1 4.575 1 4.575 1.24 4.335 1.24 4.335 1.96 6.015 1.96 6.015 1.32 6.635 1.32 6.635 0.64 6.905 0.64 6.905 0.76 6.755 0.76 6.755 1.44 6.135 1.44 6.135 2.02 6.745 2.02 6.745 1.93 6.985 1.93 ;
      POLYGON 6.275 1.16 6.035 1.16 6.035 0.54 5.675 0.54 5.675 0.62 5.655 0.62 5.655 1.56 5.535 1.56 5.535 0.62 4.935 0.62 4.935 0.54 3.855 0.54 3.855 0.62 3.235 0.62 3.235 0.6 0.835 0.6 0.835 0.66 0.255 0.66 0.255 1.39 0.315 1.39 0.315 1.63 0.195 1.63 0.195 1.51 0.135 1.51 0.135 0.54 0.715 0.54 0.715 0.48 3.355 0.48 3.355 0.5 3.735 0.5 3.735 0.42 3.935 0.42 3.935 0.4 4.175 0.4 4.175 0.42 5.055 0.42 5.055 0.5 5.555 0.5 5.555 0.42 6.155 0.42 6.155 1.04 6.275 1.04 ;
      POLYGON 5.915 1.2 5.895 1.2 5.895 1.84 5.655 1.84 5.655 1.8 5.295 1.8 5.295 1.5 4.935 1.5 4.935 1.38 5.415 1.38 5.415 1.68 5.775 1.68 5.775 1.08 5.795 1.08 5.795 0.66 5.915 0.66 ;
      POLYGON 5.315 1.22 5.195 1.22 5.195 1.1 4.815 1.1 4.815 1.84 4.455 1.84 4.455 1.72 4.695 1.72 4.695 0.66 4.815 0.66 4.815 0.98 5.315 0.98 ;
      POLYGON 4.455 0.84 4.095 0.84 4.095 1.2 3.795 1.2 3.795 1.68 3.975 1.68 3.975 1.72 4.095 1.72 4.095 1.84 3.855 1.84 3.855 1.8 3.675 1.8 3.675 1.46 3.075 1.46 3.075 1.2 3.195 1.2 3.195 1.34 3.675 1.34 3.675 1.08 3.975 1.08 3.975 0.72 4.455 0.72 ;
      POLYGON 3.555 1.22 3.435 1.22 3.435 1.08 2.955 1.08 2.955 2.04 2.835 2.04 2.835 1.08 2.395 1.08 2.395 1.16 2.155 1.16 2.155 0.96 2.835 0.96 2.835 0.72 3.115 0.72 3.115 0.84 2.955 0.84 2.955 0.96 3.555 0.96 ;
  END
END SDFFQX4

MACRO SDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFXL 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1.41 2.15 1.54 ;
        RECT 1.755 1.51 2.015 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.03 1.02 7.15 1.26 ;
        RECT 6.74 1.02 7.15 1.14 ;
        RECT 6.74 0.885 6.89 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.425 1.21 8.685 1.445 ;
        RECT 8.305 1.21 8.685 1.42 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.05 0.94 8.81 1.06 ;
        RECT 8.69 0.82 8.81 1.06 ;
        RECT 8.05 0.94 8.395 1.09 ;
        RECT 7.51 1.24 8.17 1.36 ;
        RECT 8.05 0.82 8.17 1.36 ;
        RECT 7.51 1.24 7.63 1.48 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 1.175 0.255 1.435 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.41 1.32 1.53 1.91 ;
        RECT 1.37 0.68 1.49 0.96 ;
        RECT 1.33 0.84 1.45 1.44 ;
        RECT 1.23 0.885 1.45 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
        RECT 8.53 -0.18 8.65 0.7 ;
        RECT 7.25 -0.18 7.37 0.7 ;
        RECT 5.08 0.45 5.32 0.57 ;
        RECT 5.2 -0.18 5.32 0.57 ;
        RECT 3.2 0.67 3.44 0.79 ;
        RECT 3.24 -0.18 3.36 0.79 ;
        RECT 1.79 -0.18 1.91 0.4 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
        RECT 8.53 1.92 8.65 2.79 ;
        RECT 7.09 1.92 7.21 2.79 ;
        RECT 5.04 2.23 5.16 2.79 ;
        RECT 3.38 2.17 3.62 2.29 ;
        RECT 3.38 2.17 3.5 2.79 ;
        RECT 1.83 1.79 1.95 2.79 ;
        RECT 0.555 1.46 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.07 2.04 8.95 2.04 8.95 1.685 8.09 1.685 8.09 1.66 7.97 1.66 7.97 1.54 8.21 1.54 8.21 1.565 8.95 1.565 8.95 0.46 9.07 0.46 ;
      POLYGON 8.01 0.7 7.93 0.7 7.93 1.12 7.39 1.12 7.39 1.6 7.45 1.6 7.45 1.72 7.85 1.72 7.85 2.04 7.73 2.04 7.73 1.84 7.33 1.84 7.33 1.72 6.54 1.72 6.54 1.81 6.22 1.81 6.22 1.69 6.42 1.69 6.42 0.82 6.38 0.82 6.38 0.7 6.62 0.7 6.62 0.82 6.54 0.82 6.54 1.6 7.27 1.6 7.27 1 7.81 1 7.81 0.58 7.89 0.58 7.89 0.46 8.01 0.46 ;
      POLYGON 6.95 0.7 6.83 0.7 6.83 0.58 6.26 0.58 6.26 1.06 6.1 1.06 6.1 1.35 6.3 1.35 6.3 1.47 6.1 1.47 6.1 1.93 6.85 1.93 6.85 2.05 5.98 2.05 5.98 0.94 6.14 0.94 6.14 0.58 5.56 0.58 5.56 0.81 4.84 0.81 4.84 0.52 4.48 0.52 4.48 1.17 4.6 1.17 4.6 1.29 4.36 1.29 4.36 0.4 4.96 0.4 4.96 0.69 5.44 0.69 5.44 0.46 5.62 0.46 5.62 0.36 5.86 0.36 5.86 0.46 6.95 0.46 ;
      POLYGON 6.02 0.82 5.86 0.82 5.86 1.87 5.74 1.87 5.74 1.41 4.96 1.41 4.96 1.29 5.74 1.29 5.74 0.7 6.02 0.7 ;
      POLYGON 5.78 2.25 5.43 2.25 5.43 2.11 4.6 2.11 4.6 2.25 4.36 2.25 4.36 2.11 3.84 2.11 3.84 2.05 2.515 2.05 2.515 2.03 2.25 2.03 2.25 1.67 2.27 1.67 2.27 0.74 2.51 0.74 2.51 0.86 2.39 0.86 2.39 1.79 2.37 1.79 2.37 1.91 2.635 1.91 2.635 1.93 3.84 1.93 3.84 1.27 3.76 1.27 3.76 1.15 4 1.15 4 1.27 3.96 1.27 3.96 1.99 5.55 1.99 5.55 2.13 5.78 2.13 ;
      POLYGON 5.52 1.17 4.84 1.17 4.84 1.75 4.68 1.75 4.68 1.87 4.56 1.87 4.56 1.63 4.72 1.63 4.72 1.05 4.6 1.05 4.6 0.64 4.72 0.64 4.72 0.93 4.84 0.93 4.84 1.05 5.52 1.05 ;
      POLYGON 4.32 1.81 4.08 1.81 4.08 1.69 4.12 1.69 4.12 0.88 3.875 0.88 3.875 1.03 2.96 1.03 2.96 0.48 2.88 0.48 2.88 0.36 3.12 0.36 3.12 0.48 3.08 0.48 3.08 0.91 3.755 0.91 3.755 0.76 4.12 0.76 4.12 0.64 4.24 0.64 4.24 1.69 4.32 1.69 ;
      POLYGON 3.64 1.39 3.02 1.39 3.02 1.69 3.14 1.69 3.14 1.81 2.9 1.81 2.9 1.27 2.72 1.27 2.72 0.72 2.63 0.72 2.63 0.62 2.15 0.62 2.15 1.2 1.57 1.2 1.57 1.08 2.03 1.08 2.03 0.5 2.75 0.5 2.75 0.6 2.84 0.6 2.84 1.15 3.02 1.15 3.02 1.27 3.64 1.27 ;
      POLYGON 1.1 0.92 1.095 0.92 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.8 0.98 0.8 0.98 0.68 1.1 0.68 ;
  END
END SDFFXL

MACRO CLKBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX20 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.54 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.02 1.26 8.62 1.38 ;
        RECT 8.135 1.23 8.395 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.6387 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.96 1.425 7.08 2.21 ;
        RECT 0.36 0.945 7.08 1.065 ;
        RECT 6.96 0.4 7.08 1.065 ;
        RECT 0.24 1.425 7.08 1.545 ;
        RECT 6.12 1.425 6.24 2.21 ;
        RECT 6.12 0.4 6.24 1.065 ;
        RECT 5.28 1.425 5.4 2.21 ;
        RECT 5.22 0.4 5.34 1.065 ;
        RECT 4.44 1.425 4.56 2.21 ;
        RECT 4.38 0.4 4.5 1.065 ;
        RECT 3.6 1.425 3.72 2.21 ;
        RECT 3.54 0.4 3.66 1.065 ;
        RECT 2.76 1.425 2.88 2.21 ;
        RECT 2.7 0.4 2.82 1.065 ;
        RECT 1.92 1.425 2.04 2.21 ;
        RECT 1.86 0.4 1.98 1.065 ;
        RECT 1.08 1.425 1.2 2.21 ;
        RECT 1.02 0.4 1.14 1.065 ;
        RECT 0.36 0.945 0.51 1.545 ;
        RECT 0.36 0.785 0.48 1.545 ;
        RECT 0.24 1.425 0.36 2.21 ;
        RECT 0.18 0.785 0.48 0.905 ;
        RECT 0.18 0.4 0.3 0.905 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.06 -0.18 9.18 0.72 ;
        RECT 8.22 -0.18 8.34 0.72 ;
        RECT 7.38 -0.18 7.5 0.91 ;
        RECT 6.54 -0.18 6.66 0.825 ;
        RECT 5.64 -0.18 5.76 0.825 ;
        RECT 4.8 -0.18 4.92 0.825 ;
        RECT 3.96 -0.18 4.08 0.825 ;
        RECT 3.12 -0.18 3.24 0.825 ;
        RECT 2.28 -0.18 2.4 0.825 ;
        RECT 1.44 -0.18 1.56 0.825 ;
        RECT 0.6 -0.18 0.72 0.825 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.06 1.74 9.18 2.79 ;
        RECT 8.22 1.74 8.34 2.79 ;
        RECT 7.38 1.56 7.5 2.79 ;
        RECT 6.54 1.665 6.66 2.79 ;
        RECT 5.7 1.665 5.82 2.79 ;
        RECT 4.86 1.665 4.98 2.79 ;
        RECT 4.02 1.665 4.14 2.79 ;
        RECT 3.18 1.665 3.3 2.79 ;
        RECT 2.34 1.665 2.46 2.79 ;
        RECT 1.5 1.665 1.62 2.79 ;
        RECT 0.66 1.665 0.78 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.6 0.96 7.9 0.96 7.9 1.5 9.6 1.5 9.6 2.21 9.48 2.21 9.48 1.62 8.76 1.62 8.76 2.21 8.64 2.21 8.64 1.62 7.92 1.62 7.92 2.21 7.8 2.21 7.8 1.62 7.78 1.62 7.78 1.305 0.82 1.305 0.82 1.185 7.78 1.185 7.78 0.84 7.8 0.84 7.8 0.67 7.92 0.67 7.92 0.84 8.64 0.84 8.64 0.67 8.76 0.67 8.76 0.84 9.48 0.84 9.48 0.67 9.6 0.67 ;
  END
END CLKBUFX20

MACRO OAI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X2 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.185 0.565 1.4 ;
        RECT 0.355 1.185 0.475 1.595 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.52 0.855 1.715 ;
        RECT 0.735 1.31 0.855 1.715 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.525 4.865 1.645 ;
        RECT 4.745 1.22 4.865 1.645 ;
        RECT 3.585 1.23 4.045 1.38 ;
        RECT 3.785 1.23 3.905 1.645 ;
        RECT 3.585 1.23 3.905 1.42 ;
        RECT 3.585 1.18 3.705 1.42 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 1.18 4.625 1.405 ;
        RECT 4.165 1.2 4.625 1.4 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.525 0.65 4.765 0.77 ;
        RECT 3.345 0.94 4.645 1.06 ;
        RECT 4.525 0.65 4.645 1.06 ;
        RECT 4.065 1.765 4.185 2.21 ;
        RECT 3.345 1.765 4.185 1.885 ;
        RECT 3.685 0.65 3.925 0.77 ;
        RECT 3.685 0.65 3.805 1.06 ;
        RECT 3.345 0.94 3.465 1.885 ;
        RECT 2.335 1.55 3.465 1.67 ;
        RECT 2.545 1.55 2.665 2.21 ;
        RECT 2.335 1.52 2.595 1.67 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 2.845 0.46 3.085 0.58 ;
        RECT 2.845 -0.18 2.965 0.58 ;
        RECT 2.005 0.46 2.245 0.58 ;
        RECT 2.005 -0.18 2.125 0.58 ;
        RECT 0.615 -0.18 0.735 0.825 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 4.705 1.765 4.825 2.79 ;
        RECT 3.265 2.005 3.505 2.15 ;
        RECT 3.265 2.005 3.385 2.79 ;
        RECT 1.905 1.56 2.025 2.79 ;
        RECT 0.595 1.835 0.715 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.125 0.65 5.005 0.65 5.005 0.53 4.285 0.53 4.285 0.65 4.165 0.65 4.165 0.53 3.445 0.53 3.445 0.65 3.415 0.65 3.415 0.82 1.705 0.82 1.705 0.77 1.585 0.77 1.585 0.65 1.825 0.65 1.825 0.7 2.425 0.7 2.425 0.65 2.665 0.65 2.665 0.7 3.295 0.7 3.295 0.41 5.125 0.41 ;
      POLYGON 3.225 1.4 1.215 1.4 1.215 1.52 1.135 1.52 1.135 1.955 1.015 1.955 1.015 1.4 1.095 1.4 1.095 0.6 1.215 0.6 1.215 1.28 3.225 1.28 ;
      POLYGON 2.445 1.09 1.345 1.09 1.345 0.48 0.975 0.48 0.975 1.065 0.185 1.065 0.185 1.715 0.295 1.715 0.295 1.955 0.175 1.955 0.175 1.835 0.065 1.835 0.065 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.945 0.855 0.945 0.855 0.36 1.465 0.36 1.465 0.97 2.445 0.97 ;
  END
END OAI2BB2X2

MACRO FILL32
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILL32 0 0 ;
  SIZE 9.28 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.28 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.28 0.18 ;
    END
  END VSS
END FILL32

MACRO OAI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.01 2.54 1.465 ;
        RECT 2.39 1.01 2.51 1.495 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 1.055 2.05 1.295 ;
        RECT 1.81 1.175 2.005 1.435 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.04 1.38 1.495 ;
        RECT 1.25 1.01 1.37 1.495 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.465 ;
        RECT 0.36 1.01 0.48 1.495 ;
    END
  END A0
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.57 1.02 1.69 1.435 ;
        RECT 1.52 1.095 1.67 1.495 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.15 1.09 1.435 ;
        RECT 0.83 1.02 0.95 1.295 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.466 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 1.465 2.83 1.725 ;
        RECT 1.83 0.77 2.79 0.89 ;
        RECT 2.67 0.6 2.79 0.89 ;
        RECT 1.41 1.615 2.78 1.735 ;
        RECT 2.66 0.77 2.78 1.735 ;
        RECT 1.83 0.6 1.95 0.89 ;
        RECT 1.41 1.615 1.53 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 0.99 -0.18 1.11 0.65 ;
        RECT 0.15 -0.18 0.27 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.37 1.855 2.49 2.79 ;
        RECT 0.35 1.615 0.47 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.37 0.65 2.25 0.65 2.25 0.53 2.07 0.53 2.07 0.48 1.53 0.48 1.53 0.89 0.57 0.89 0.57 0.6 0.69 0.6 0.69 0.77 1.41 0.77 1.41 0.36 2.19 0.36 2.19 0.41 2.37 0.41 ;
  END
END OAI33X1

MACRO SDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX4 0 0 ;
  SIZE 13.34 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 1.1 0.525 1.34 ;
        RECT 0.07 1.175 0.525 1.295 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.09 1.04 1.21 1.43 ;
        RECT 0.885 1.19 1.21 1.41 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.2 1.725 1.41 ;
        RECT 1.605 1.04 1.725 1.41 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.175 3.41 1.435 ;
        RECT 3.12 1.175 3.41 1.295 ;
        RECT 3.12 1.055 3.24 1.295 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 1.175 3.7 1.535 ;
        RECT 3.53 1 3.65 1.365 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.185 0.72 10.385 0.84 ;
        RECT 10.245 1.44 10.365 2.21 ;
        RECT 10.065 1.44 10.365 1.56 ;
        RECT 9.38 1.32 10.185 1.44 ;
        RECT 9.405 0.72 9.525 2.21 ;
        RECT 9.35 1.175 9.525 1.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.105 0.72 12.305 0.84 ;
        RECT 11.925 1.32 12.045 2.21 ;
        RECT 11.09 1.32 12.045 1.44 ;
        RECT 11.12 0.72 11.24 1.56 ;
        RECT 11.085 1.44 11.205 2.21 ;
        RECT 11.09 1.175 11.24 1.56 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.34 0.18 ;
        RECT 12.665 -0.18 12.785 0.71 ;
        RECT 11.585 -0.18 11.825 0.36 ;
        RECT 10.625 -0.18 10.865 0.36 ;
        RECT 9.665 -0.18 9.905 0.36 ;
        RECT 8.705 -0.18 8.945 0.36 ;
        RECT 7.865 -0.18 7.985 0.9 ;
        RECT 6.145 -0.18 6.385 0.32 ;
        RECT 4.215 -0.18 4.335 0.92 ;
        RECT 3.22 -0.18 3.34 0.88 ;
        RECT 1.23 -0.18 1.35 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.34 2.79 ;
        RECT 12.345 1.58 12.465 2.79 ;
        RECT 11.505 1.56 11.625 2.79 ;
        RECT 10.665 1.56 10.785 2.79 ;
        RECT 9.825 1.56 9.945 2.79 ;
        RECT 8.985 1.56 9.105 2.79 ;
        RECT 8.085 1.62 8.205 2.79 ;
        RECT 6.205 1.74 6.325 2.79 ;
        RECT 4.3 1.98 4.42 2.79 ;
        RECT 3.22 1.94 3.34 2.79 ;
        RECT 1.29 2.01 1.41 2.79 ;
        RECT 0.39 1.59 0.51 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.205 0.9 13.025 0.9 13.025 1.46 12.885 1.46 12.885 2.21 12.765 2.21 12.765 1.46 12.165 1.46 12.165 1.3 12.405 1.3 12.405 1.34 12.905 1.34 12.905 0.78 13.085 0.78 13.085 0.66 13.205 0.66 ;
      POLYGON 12.745 1.22 12.625 1.22 12.625 0.95 12.425 0.95 12.425 0.6 8.935 0.6 8.935 0.66 8.405 0.66 8.405 0.78 8.765 0.78 8.765 1.28 9.23 1.28 9.23 1.4 8.625 1.4 8.625 2.14 8.505 2.14 8.505 1.4 8.125 1.4 8.125 1.5 8.005 1.5 8.005 1.26 8.125 1.26 8.125 1.28 8.645 1.28 8.645 0.9 8.285 0.9 8.285 0.54 8.815 0.54 8.815 0.48 12.545 0.48 12.545 0.83 12.745 0.83 ;
      POLYGON 8.525 1.16 8.285 1.16 8.285 1.14 7.885 1.14 7.885 1.76 7.545 1.76 7.545 1.8 7.305 1.8 7.305 1.68 7.425 1.68 7.425 1.64 7.765 1.64 7.765 1.14 7.225 1.14 7.225 0.66 7.345 0.66 7.345 1.02 8.525 1.02 ;
      POLYGON 7.645 1.52 7.525 1.52 7.525 1.38 6.985 1.38 6.985 0.54 6.625 0.54 6.625 0.56 5.905 0.56 5.905 0.54 5.385 0.54 5.385 1.36 5.445 1.36 5.445 1.48 5.205 1.48 5.205 1.36 5.265 1.36 5.265 0.54 4.855 0.54 4.855 0.68 4.755 0.68 4.755 0.8 4.845 0.8 4.845 1.58 4.725 1.58 4.725 0.92 4.635 0.92 4.635 0.56 4.735 0.56 4.735 0.42 5.665 0.42 5.665 0.38 5.905 0.38 5.905 0.42 6.025 0.42 6.025 0.44 6.505 0.44 6.505 0.42 7.105 0.42 7.105 1.26 7.645 1.26 ;
      POLYGON 6.865 1.86 6.745 1.86 6.745 1.48 6.005 1.48 6.005 1.36 6.745 1.36 6.745 0.66 6.865 0.66 ;
      POLYGON 6.625 1.24 5.685 1.24 5.685 1.86 5.565 1.86 5.565 0.84 5.505 0.84 5.505 0.72 5.745 0.72 5.745 0.84 5.685 0.84 5.685 1.12 6.625 1.12 ;
      POLYGON 5.245 1.86 4.18 1.86 4.18 2.24 3.46 2.24 3.46 1.82 2.965 1.82 2.965 1.94 2.7 1.94 2.7 2.06 2.58 2.06 2.58 1.94 2.44 1.94 2.44 0.7 2.76 0.7 2.76 0.82 2.56 0.82 2.56 1.82 2.845 1.82 2.845 1.7 3.58 1.7 3.58 2.12 4.06 2.12 4.06 1.74 4.965 1.74 4.965 1.12 5.025 1.12 5.025 0.66 5.145 0.66 5.145 1.24 5.085 1.24 5.085 1.62 5.245 1.62 ;
      POLYGON 4.605 1.18 3.94 1.18 3.94 2 3.7 2 3.7 1.88 3.82 1.88 3.82 0.88 3.64 0.88 3.64 0.64 3.76 0.64 3.76 0.76 3.94 0.76 3.94 1.06 4.605 1.06 ;
      POLYGON 3 1.58 2.68 1.58 2.68 1.46 2.88 1.46 2.88 0.52 1.805 0.52 1.805 0.68 1.77 0.68 1.77 0.8 1.965 0.8 1.965 1.65 1.71 1.65 1.71 1.53 1.845 1.53 1.845 0.92 1.65 0.92 1.65 0.56 1.685 0.56 1.685 0.4 2.36 0.4 2.36 0.36 2.6 0.36 2.6 0.4 3 0.4 ;
      POLYGON 2.28 2.06 2.16 2.06 2.16 1.89 0.81 1.89 0.81 1.65 0.645 1.65 0.645 0.86 0.53 0.86 0.53 0.74 0.77 0.74 0.77 0.86 0.765 0.86 0.765 1.53 0.93 1.53 0.93 1.77 2.16 1.77 2.16 0.64 2.28 0.64 ;
  END
END SDFFTRX4

MACRO NOR2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BXL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1 0.51 1.49 ;
        RECT 0.36 1 0.51 1.465 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.235 1.36 ;
        RECT 1.115 1.12 1.235 1.36 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.12 0.76 0.675 0.88 ;
        RECT 0.555 0.4 0.675 0.88 ;
        RECT 0.335 1.61 0.455 1.85 ;
        RECT 0.12 1.61 0.455 1.73 ;
        RECT 0.07 1.465 0.24 1.725 ;
        RECT 0.12 0.76 0.24 1.73 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.975 -0.18 1.095 0.64 ;
        RECT 0.135 -0.18 0.255 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.975 1.61 1.095 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.73 1.395 1.73 1.395 1 0.815 1 0.815 0.76 0.935 0.76 0.935 0.88 1.395 0.88 1.395 0.4 1.515 0.4 ;
  END
END NOR2BXL

MACRO MXI2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.76 0.51 1.21 ;
        RECT 0.36 0.76 0.48 1.37 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.23 1.8 1.445 ;
        RECT 1.465 1.23 1.725 1.465 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.99 2.12 1.11 ;
        RECT 1.22 0.97 2.015 1.09 ;
        RECT 1.755 0.94 2.015 1.11 ;
        RECT 1.44 0.41 1.56 1.09 ;
        RECT 0.7 0.41 1.56 0.53 ;
        RECT 0.7 0.41 0.82 1.43 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.65 1.32 0.77 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.94 0.65 1.06 1.67 ;
        RECT 0.93 1.55 1.05 2.2 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.78 -0.18 1.9 0.82 ;
        RECT 0.2 -0.18 0.32 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.71 1.825 1.83 2.79 ;
        RECT 0.2 1.55 0.32 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.36 1.825 2.25 1.825 2.25 2.065 2.13 2.065 2.13 1.705 1.21 1.705 1.21 1.23 1.33 1.23 1.33 1.585 2.24 1.585 2.24 0.82 2.2 0.82 2.2 0.58 2.32 0.58 2.32 0.7 2.36 0.7 ;
  END
END MXI2X1

MACRO NOR4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 1.02 0.365 1.26 ;
        RECT 0.07 1.02 0.365 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 1.25 2.89 1.5 ;
        RECT 2.625 1.23 2.885 1.5 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.52 1.34 1.64 1.725 ;
        RECT 1.43 1.22 1.55 1.46 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.995 1.22 1.115 1.46 ;
        RECT 0.94 1.465 1.09 1.725 ;
        RECT 0.97 1.34 1.09 1.725 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4572 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.07 1.465 2.25 1.725 ;
        RECT 1.315 0.71 2.215 0.83 ;
        RECT 2.095 0.59 2.215 0.83 ;
        RECT 0.95 1.845 2.19 1.965 ;
        RECT 2.07 0.71 2.19 1.965 ;
        RECT 1.195 0.65 1.435 0.77 ;
        RECT 0.95 1.845 1.07 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.515 -0.18 2.635 0.83 ;
        RECT 1.615 0.46 1.855 0.58 ;
        RECT 1.615 -0.18 1.735 0.58 ;
        RECT 0.775 -0.18 0.895 0.53 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.31 1.845 2.43 2.79 ;
        RECT 0.135 1.98 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.13 1.74 2.97 1.74 2.97 1.86 2.85 1.86 2.85 1.62 3.01 1.62 3.01 1.11 2.31 1.11 2.31 0.99 2.935 0.99 2.935 0.59 3.055 0.59 3.055 0.87 3.13 0.87 ;
      POLYGON 1.95 1.1 0.68 1.1 0.68 1.58 0.56 1.58 0.56 0.98 0.525 0.98 0.525 0.68 0.645 0.68 0.645 0.86 0.68 0.86 0.68 0.98 1.95 0.98 ;
  END
END NOR4BBX1

MACRO CLKINVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX2 0 0 ;
  SIZE 1.45 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 1 0.49 1.24 ;
        RECT 0.07 1.025 0.49 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.885 0.8 1.145 ;
        RECT 0.65 0.68 0.77 2.01 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.45 0.18 ;
        RECT 1.07 -0.18 1.19 0.73 ;
        RECT 0.23 -0.18 0.35 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.45 2.79 ;
        RECT 1.07 1.36 1.19 2.79 ;
        RECT 0.23 1.36 0.35 2.79 ;
    END
  END VDD
END CLKINVX2

MACRO SDFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX2 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 1.09 1.38 1.59 ;
        RECT 1.23 1.09 1.38 1.56 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.87 1.19 6.18 1.43 ;
        RECT 5.87 1.175 6.02 1.435 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 1.21 7.815 1.41 ;
        RECT 7.34 1.21 7.815 1.38 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.74 0.97 7.9 1.09 ;
        RECT 7.08 0.94 7.525 1.09 ;
        RECT 7.08 0.91 7.2 1.15 ;
        RECT 6.54 1.23 6.86 1.35 ;
        RECT 6.74 0.97 6.86 1.35 ;
        RECT 6.54 1.23 6.66 1.47 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.68 0.72 2.04 ;
        RECT 0.36 0.885 0.72 1.145 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 7.56 -0.18 7.68 0.79 ;
        RECT 6.26 -0.18 6.38 0.79 ;
        RECT 4.13 -0.18 4.37 0.37 ;
        RECT 2.25 0.63 2.49 0.75 ;
        RECT 2.25 -0.18 2.37 0.75 ;
        RECT 1.02 -0.18 1.14 0.73 ;
        RECT 0.18 -0.18 0.3 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.44 1.91 7.56 2.79 ;
        RECT 6.16 1.91 6.28 2.79 ;
        RECT 4.11 2.23 4.23 2.79 ;
        RECT 2.27 2.01 2.51 2.13 ;
        RECT 2.27 2.01 2.39 2.79 ;
        RECT 1.02 1.68 1.14 2.79 ;
        RECT 0.18 1.39 0.3 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.14 1.77 7.98 1.77 7.98 2.03 7.86 2.03 7.86 1.65 7.1 1.65 7.1 1.43 6.98 1.43 6.98 1.31 7.22 1.31 7.22 1.53 8.02 1.53 8.02 0.79 7.98 0.79 7.98 0.55 8.1 0.55 8.1 0.67 8.14 0.67 ;
      POLYGON 7.04 0.79 6.62 0.79 6.62 1.11 6.42 1.11 6.42 1.59 6.92 1.59 6.92 2.03 6.8 2.03 6.8 1.71 5.61 1.71 5.61 1.81 5.29 1.81 5.29 1.69 5.49 1.69 5.49 0.91 5.43 0.91 5.43 0.67 5.55 0.67 5.55 0.79 5.61 0.79 5.61 1.59 6.3 1.59 6.3 0.99 6.5 0.99 6.5 0.67 6.92 0.67 6.92 0.55 7.04 0.55 ;
      POLYGON 5.96 0.79 5.84 0.79 5.84 0.55 5.31 0.55 5.31 1.09 5.17 1.09 5.17 1.37 5.37 1.37 5.37 1.49 5.17 1.49 5.17 1.93 5.92 1.93 5.92 2.05 5.05 2.05 5.05 0.97 5.19 0.97 5.19 0.55 4.61 0.55 4.61 0.61 3.53 0.61 3.53 1.23 3.41 1.23 3.41 0.49 4.49 0.49 4.49 0.43 4.69 0.43 4.69 0.41 4.93 0.41 4.93 0.43 5.96 0.43 ;
      POLYGON 5.07 0.85 4.93 0.85 4.93 1.87 4.81 1.87 4.81 1.49 3.89 1.49 3.89 1.37 4.81 1.37 4.81 0.73 5.07 0.73 ;
      POLYGON 4.85 2.25 4.35 2.25 4.35 2.11 3.53 2.11 3.53 2.25 3.29 2.25 3.29 2.11 2.83 2.11 2.83 1.89 1.56 1.89 1.56 1.95 1.44 1.95 1.44 1.71 1.5 1.71 1.5 0.68 1.62 0.68 1.62 1.77 2.83 1.77 2.83 1.23 2.81 1.23 2.81 1.11 3.05 1.11 3.05 1.23 2.95 1.23 2.95 1.99 4.47 1.99 4.47 2.13 4.85 2.13 ;
      POLYGON 4.49 1.25 3.77 1.25 3.77 1.75 3.75 1.75 3.75 1.87 3.63 1.87 3.63 1.63 3.65 1.63 3.65 0.73 3.89 0.73 3.89 0.85 3.77 0.85 3.77 1.13 4.49 1.13 ;
      POLYGON 3.33 1.87 3.21 1.87 3.21 1.47 3.17 1.47 3.17 0.91 2.82 0.91 2.82 0.99 2.29 0.99 2.29 1.23 2.17 1.23 2.17 0.87 2.7 0.87 2.7 0.79 3.13 0.79 3.13 0.67 3.25 0.67 3.25 0.79 3.29 0.79 3.29 1.35 3.33 1.35 ;
      POLYGON 2.71 1.47 2.03 1.47 2.03 1.65 1.79 1.65 1.79 1.53 1.91 1.53 1.91 0.91 1.89 0.91 1.89 0.67 1.79 0.67 1.79 0.56 1.38 0.56 1.38 0.97 1 0.97 1 1.24 0.88 1.24 0.88 0.85 1.26 0.85 1.26 0.44 1.91 0.44 1.91 0.55 2.01 0.55 2.01 0.79 2.03 0.79 2.03 1.35 2.71 1.35 ;
  END
END SDFFQX2

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.735 0.82 1.17 ;
        RECT 0.65 0.595 0.8 1.005 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.21 0.795 1.38 1.215 ;
        RECT 1.21 0.795 1.33 1.235 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.785 1.67 1.235 ;
        RECT 1.53 0.76 1.65 1.235 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.885 0.51 1.34 ;
        RECT 0.38 0.885 0.5 1.36 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3478 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.355 1.515 2.01 ;
        RECT 0.97 1.355 1.515 1.475 ;
        RECT 0.94 1.175 1.09 1.435 ;
        RECT 0.97 0.59 1.09 1.475 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.69 -0.18 1.81 0.64 ;
        RECT 0.22 -0.18 0.34 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 0.555 1.835 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 2.25 0.975 2.25 0.975 1.715 0.255 1.715 0.255 2.21 0.135 2.21 0.135 1.56 0.255 1.56 0.255 1.595 1.095 1.595 1.095 2.13 1.815 2.13 1.815 1.56 1.935 1.56 ;
  END
END AOI22X1

MACRO AO21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.4 1.67 1.735 ;
        RECT 1.4 1.355 1.64 1.52 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.2 1.17 1.32 ;
        RECT 1.05 1.08 1.17 1.32 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.065 0.53 1.5 ;
        RECT 0.41 1.04 0.53 1.5 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 1.4 2.825 1.52 ;
        RECT 2.13 0.68 2.25 1.52 ;
        RECT 2.1 0.885 2.25 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.65 0.74 1.89 0.86 ;
        RECT 1.65 -0.18 1.77 0.86 ;
        RECT 0.55 -0.18 0.67 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.18 1.98 2.3 2.79 ;
        RECT 0.8 1.86 0.92 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.97 1.24 1.91 1.24 1.91 1.98 1.79 1.98 1.79 1.1 1.29 1.1 1.29 0.68 1.41 0.68 1.41 0.98 1.91 0.98 1.91 1 1.97 1 ;
      POLYGON 1.4 1.92 1.16 1.92 1.16 1.74 0.56 1.74 0.56 1.92 0.32 1.92 0.32 1.8 0.44 1.8 0.44 1.62 1.28 1.62 1.28 1.8 1.4 1.8 ;
  END
END AO21XL

MACRO OAI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32XL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.175 2.54 1.435 ;
        RECT 2.165 1.175 2.54 1.295 ;
        RECT 2.165 1.055 2.285 1.295 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.36 1.295 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1.465 2.25 1.725 ;
        RECT 1.845 1.535 2.25 1.655 ;
        RECT 1.845 1.415 1.965 1.655 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.175 0.82 1.61 ;
        RECT 0.65 1.175 0.82 1.59 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.34 0.51 1.755 ;
        RECT 0.36 1.03 0.48 1.755 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 1.175 2 1.295 ;
        RECT 1.88 0.635 2 1.295 ;
        RECT 1.465 1.52 1.725 1.67 ;
        RECT 1.585 1.175 1.705 1.995 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 0.98 0.695 1.22 0.815 ;
        RECT 0.98 -0.18 1.1 0.815 ;
        RECT 0.2 -0.18 0.32 0.875 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 2.325 1.875 2.445 2.79 ;
        RECT 0.2 1.875 0.32 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.42 0.875 2.3 0.875 2.3 0.515 1.58 0.515 1.58 1.055 0.62 1.055 0.62 0.635 0.74 0.635 0.74 0.935 1.46 0.935 1.46 0.395 2.42 0.395 ;
  END
END OAI32XL

MACRO NOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 1.28 0.82 1.755 ;
        RECT 0.65 1.28 0.82 1.73 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.35 1.34 0.53 1.725 ;
        RECT 0.36 1.33 0.51 1.725 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 1.28 1.17 1.65 ;
        RECT 0.94 1.36 1.09 1.725 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 1.04 1.53 1.16 ;
        RECT 1.41 0.68 1.53 1.16 ;
        RECT 1.29 0.885 1.41 1.89 ;
        RECT 1.21 1.77 1.33 2.01 ;
        RECT 1.23 0.885 1.53 1.16 ;
        RECT 0.57 0.68 0.69 1.16 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 0.99 -0.18 1.11 0.92 ;
        RECT 0.135 -0.18 0.255 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.22 1.845 0.34 2.79 ;
    END
  END VDD
END NOR3XL

MACRO AOI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X2 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.205 0.94 3.525 1.16 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.625 0.94 2.885 1.155 ;
        RECT 2.505 0.94 2.885 1.13 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.555 0.99 1.795 1.11 ;
        RECT 0.595 0.94 1.675 1.06 ;
        RECT 0.435 0.99 0.855 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.055 1.18 1.435 1.4 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6208 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.385 1.28 3.505 1.99 ;
        RECT 2.265 1.28 3.505 1.4 ;
        RECT 3.125 0.65 3.365 0.77 ;
        RECT 1.195 0.7 3.245 0.82 ;
        RECT 2.265 0.65 2.505 0.82 ;
        RECT 2.265 0.65 2.385 1.4 ;
        RECT 2.1 0.7 2.385 1.145 ;
        RECT 1.075 0.65 1.315 0.77 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.605 -0.18 3.725 0.64 ;
        RECT 2.685 0.46 2.925 0.58 ;
        RECT 2.685 -0.18 2.805 0.58 ;
        RECT 1.845 0.46 2.085 0.58 ;
        RECT 1.845 -0.18 1.965 0.58 ;
        RECT 0.335 -0.18 0.455 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 1.875 2.14 1.995 2.79 ;
        RECT 0.975 1.76 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.925 2.23 2.185 2.23 2.185 1.88 2.065 1.88 2.065 1.76 2.305 1.76 2.305 2.11 2.965 2.11 2.965 1.52 3.085 1.52 3.085 2.11 3.805 2.11 3.805 1.34 3.925 1.34 ;
      POLYGON 2.665 1.99 2.545 1.99 2.545 1.64 1.515 1.64 1.515 2.21 1.395 2.21 1.395 1.64 0.675 1.64 0.675 2.21 0.555 2.21 0.555 1.52 2.665 1.52 ;
  END
END AOI211X2

MACRO MX4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X2 0 0 ;
  SIZE 7.25 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.79 0.885 1.96 1.155 ;
        RECT 1.73 1.035 1.87 1.285 ;
    END
  END S1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.95 1.08 3.07 1.32 ;
        RECT 2.68 1.175 3.07 1.295 ;
        RECT 2.68 1.175 2.83 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.13 1.4 4.3 1.835 ;
        RECT 4.17 1.38 4.3 1.835 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.49 1.38 4.67 1.63 ;
        RECT 4.42 1.46 4.625 1.725 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.05 1.2 6.365 1.415 ;
        RECT 6.05 1.2 6.17 1.56 ;
    END
  END D
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2976 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.6533 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.485 1.175 6.89 1.435 ;
        RECT 6.485 0.96 6.605 1.435 ;
        RECT 5.71 0.96 6.605 1.08 ;
        RECT 5.71 0.96 5.83 1.22 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.35 1.57 2.59 1.69 ;
        RECT 2.47 0.66 2.59 1.025 ;
        RECT 2.42 0.885 2.54 1.69 ;
        RECT 2.39 0.885 2.54 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.25 0.18 ;
        RECT 6.15 0.72 6.39 0.84 ;
        RECT 6.15 -0.18 6.27 0.84 ;
        RECT 4.45 0.54 4.69 0.66 ;
        RECT 4.57 -0.18 4.69 0.66 ;
        RECT 2.95 -0.18 3.07 0.38 ;
        RECT 1.99 -0.18 2.11 0.525 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.25 2.79 ;
        RECT 6.21 1.92 6.33 2.79 ;
        RECT 4.34 2.195 4.58 2.79 ;
        RECT 2.83 2.05 3.07 2.17 ;
        RECT 2.83 2.05 2.95 2.79 ;
        RECT 1.87 2.29 2.11 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.13 1.92 6.75 1.92 6.75 2.04 6.63 2.04 6.63 1.8 5.91 1.8 5.91 2.22 5.19 2.22 5.19 2.075 3.89 2.075 3.89 1.74 3.84 1.74 3.84 1.48 3.96 1.48 3.96 1.62 4.01 1.62 4.01 1.955 5.19 1.955 5.19 1 5.31 1 5.31 2.1 5.79 2.1 5.79 1.74 5.73 1.74 5.73 1.46 5.85 1.46 5.85 1.62 5.91 1.62 5.91 1.68 7.01 1.68 7.01 1.055 6.725 1.055 6.725 0.66 6.845 0.66 6.845 0.935 7.13 0.935 ;
      POLYGON 5.67 1.98 5.43 1.98 5.43 0.88 4.965 0.88 4.965 0.9 4.05 0.9 4.05 0.54 3.375 0.54 3.375 0.62 2.71 0.62 2.71 0.54 2.35 0.54 2.35 0.765 1.75 0.765 1.75 0.49 1.215 0.49 1.215 0.93 1.24 0.93 1.24 1.65 1.18 1.65 1.18 1.77 1.06 1.77 1.06 1.53 1.12 1.53 1.12 1.05 1.095 1.05 1.095 0.37 1.87 0.37 1.87 0.645 2.23 0.645 2.23 0.42 2.83 0.42 2.83 0.5 3.255 0.5 3.255 0.42 4.17 0.42 4.17 0.78 4.845 0.78 4.845 0.76 5.43 0.76 5.43 0.66 5.55 0.66 5.55 1.86 5.67 1.86 ;
      POLYGON 5.03 1.42 4.79 1.42 4.79 1.26 3.72 1.26 3.72 1.58 3.55 1.58 3.55 1.7 3.43 1.7 3.43 1.46 3.6 1.46 3.6 1.14 3.97 1.14 3.97 1.02 4.09 1.02 4.09 1.14 5.03 1.14 ;
      POLYGON 3.93 0.9 3.48 0.9 3.48 1.34 3.31 1.34 3.31 1.82 3.65 1.82 3.65 1.86 3.77 1.86 3.77 1.98 3.53 1.98 3.53 1.94 3.19 1.94 3.19 1.93 2.25 1.93 2.25 2.17 1.665 2.17 1.665 2.25 0.22 2.25 0.22 1.44 0.08 1.44 0.08 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.84 0.2 0.84 0.2 1.32 0.34 1.32 0.34 2.13 1.545 2.13 1.545 2.05 2.13 2.05 2.13 1.81 3.19 1.81 3.19 1.22 3.36 1.22 3.36 0.78 3.81 0.78 3.81 0.66 3.93 0.66 ;
      POLYGON 2.27 1.41 2.23 1.41 2.23 1.53 2.01 1.53 2.01 1.93 1.425 1.93 1.425 2.01 0.64 2.01 0.64 1.64 0.615 1.64 0.615 0.6 0.735 0.6 0.735 1.52 0.76 1.52 0.76 1.89 1.305 1.89 1.305 1.81 1.89 1.81 1.89 1.41 2.11 1.41 2.11 1.29 2.15 1.29 2.15 1.17 2.27 1.17 ;
      POLYGON 1.63 0.915 1.51 0.915 1.51 1.57 1.63 1.57 1.63 1.69 1.39 1.69 1.39 1.41 1.36 1.41 1.36 1.17 1.39 1.17 1.39 0.795 1.51 0.795 1.51 0.61 1.63 0.61 ;
      POLYGON 1 1.41 0.88 1.41 0.88 1.29 0.855 1.29 0.855 0.48 0.495 0.48 0.495 1.2 0.32 1.2 0.32 0.96 0.375 0.96 0.375 0.36 0.975 0.36 0.975 1.17 1 1.17 ;
  END
END MX4X2

MACRO NAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X6 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.915 0.99 5.035 1.345 ;
        RECT 0.65 0.99 5.035 1.11 ;
        RECT 3.425 0.99 3.665 1.195 ;
        RECT 1.915 0.99 2.155 1.195 ;
        RECT 0.435 1.08 0.8 1.2 ;
        RECT 0.65 0.885 0.8 1.2 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.785 1.3 4.175 1.42 ;
        RECT 3.785 1.23 4.045 1.42 ;
        RECT 1.295 1.315 3.905 1.435 ;
        RECT 2.655 1.3 2.895 1.435 ;
        RECT 1.175 1.28 1.415 1.4 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.7541 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.555 5.275 1.675 ;
        RECT 5.155 0.75 5.275 1.675 ;
        RECT 5 1.465 5.275 1.675 ;
        RECT 0.975 0.75 5.275 0.87 ;
        RECT 5 1.465 5.15 1.725 ;
        RECT 4.755 1.555 4.875 2.21 ;
        RECT 4.135 0.4 4.255 0.87 ;
        RECT 3.915 1.555 4.035 2.21 ;
        RECT 3.075 1.555 3.195 2.21 ;
        RECT 2.855 0.4 2.975 0.87 ;
        RECT 2.235 1.555 2.355 2.21 ;
        RECT 1.395 1.555 1.515 2.21 ;
        RECT 0.975 0.4 1.095 0.87 ;
        RECT 0.555 1.555 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 3.435 0.46 3.675 0.63 ;
        RECT 3.435 -0.18 3.555 0.63 ;
        RECT 1.655 0.46 1.895 0.63 ;
        RECT 1.655 -0.18 1.775 0.63 ;
        RECT 0.335 -0.18 0.455 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 5.175 1.845 5.295 2.79 ;
        RECT 4.335 1.795 4.455 2.79 ;
        RECT 3.495 1.795 3.615 2.79 ;
        RECT 2.655 1.795 2.775 2.79 ;
        RECT 1.815 1.795 1.935 2.79 ;
        RECT 0.975 1.795 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND2X6

MACRO TLATNTSCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX20 0 0 ;
  SIZE 16.53 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.04 0.29 1.335 ;
        RECT 0.07 1.13 0.22 1.435 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.82 1.04 0.94 1.28 ;
        RECT 0.68 1.16 0.94 1.28 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 1.23 1.435 1.38 ;
        RECT 1.18 1.1 1.42 1.38 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.608 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.1 1.205 16.22 2.205 ;
        RECT 16.1 0.405 16.22 1.03 ;
        RECT 9.35 1.205 16.22 1.325 ;
        RECT 15.92 0.91 16.22 1.03 ;
        RECT 15.26 1.03 16.04 1.325 ;
        RECT 15.26 0.405 15.38 2.21 ;
        RECT 14.42 0.405 14.54 2.21 ;
        RECT 13.58 1.03 14.54 1.325 ;
        RECT 13.58 0.405 13.7 2.21 ;
        RECT 12.74 0.405 12.86 2.21 ;
        RECT 11.9 1.03 12.86 1.325 ;
        RECT 11.9 0.405 12.02 2.21 ;
        RECT 11.06 1.205 11.18 2.21 ;
        RECT 10.88 0.79 11.18 0.91 ;
        RECT 11.06 0.405 11.18 0.91 ;
        RECT 10.22 1.03 11 1.325 ;
        RECT 10.88 0.79 11 1.325 ;
        RECT 10.22 0.405 10.34 2.21 ;
        RECT 9.38 0.4 9.5 2.21 ;
        RECT 9.35 1.175 9.5 1.435 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 16.53 0.18 ;
        RECT 15.68 -0.18 15.8 0.91 ;
        RECT 14.84 -0.18 14.96 0.91 ;
        RECT 14 -0.18 14.12 0.91 ;
        RECT 13.16 -0.18 13.28 0.91 ;
        RECT 12.32 -0.18 12.44 0.91 ;
        RECT 11.48 -0.18 11.6 0.91 ;
        RECT 10.64 -0.18 10.76 0.91 ;
        RECT 9.8 -0.18 9.92 0.91 ;
        RECT 8.96 -0.18 9.08 0.87 ;
        RECT 7.64 0.46 7.88 0.58 ;
        RECT 7.64 -0.18 7.76 0.58 ;
        RECT 6.36 0.46 6.6 0.58 ;
        RECT 6.36 -0.18 6.48 0.58 ;
        RECT 5.14 -0.18 5.26 0.64 ;
        RECT 4.3 -0.18 4.42 0.64 ;
        RECT 2.97 0.47 3.21 0.59 ;
        RECT 2.97 -0.18 3.09 0.59 ;
        RECT 0.98 -0.18 1.22 0.34 ;
        RECT 0.14 -0.18 0.26 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 16.53 2.79 ;
        RECT 15.68 1.445 15.8 2.79 ;
        RECT 14.84 1.445 14.96 2.79 ;
        RECT 14 1.445 14.12 2.79 ;
        RECT 13.16 1.445 13.28 2.79 ;
        RECT 12.32 1.445 12.44 2.79 ;
        RECT 11.48 1.445 11.6 2.79 ;
        RECT 10.64 1.445 10.76 2.79 ;
        RECT 9.8 1.445 9.92 2.79 ;
        RECT 8.96 1.71 9.08 2.79 ;
        RECT 8.12 1.71 8.24 2.79 ;
        RECT 7.28 1.71 7.4 2.79 ;
        RECT 6.44 1.71 6.56 2.79 ;
        RECT 5.6 1.71 5.72 2.79 ;
        RECT 4.7 2.03 4.94 2.15 ;
        RECT 4.7 2.03 4.82 2.79 ;
        RECT 3.74 2.06 3.98 2.18 ;
        RECT 3.74 2.06 3.86 2.79 ;
        RECT 3.07 2.03 3.19 2.79 ;
        RECT 0.98 1.5 1.1 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.23 1.23 9.02 1.23 9.02 1.59 8.66 1.59 8.66 2.21 8.54 2.21 8.54 1.59 7.82 1.59 7.82 2.21 7.7 2.21 7.7 1.59 6.98 1.59 6.98 2.21 6.86 2.21 6.86 1.59 6.14 1.59 6.14 2.21 6.02 2.21 6.02 1.59 5.3 1.59 5.3 2.21 5.18 2.21 5.18 1.47 8.9 1.47 8.9 1.11 8.34 1.11 8.34 0.82 5.84 0.82 5.84 0.77 5.72 0.77 5.72 0.65 5.96 0.65 5.96 0.7 7 0.7 7 0.65 7.24 0.65 7.24 0.7 8.34 0.7 8.34 0.59 8.46 0.59 8.46 0.99 9.02 0.99 9.02 1.11 9.23 1.11 ;
      POLYGON 8.78 1.35 5.06 1.35 5.06 1.91 3.71 1.91 3.71 1.67 2.63 1.67 2.63 1.29 2.55 1.29 2.55 1.05 2.63 1.05 2.63 0.95 3.57 0.95 3.57 0.6 3.81 0.6 3.81 0.72 3.69 0.72 3.69 1.07 2.75 1.07 2.75 1.55 3.83 1.55 3.83 1.79 4.94 1.79 4.94 1.23 8.78 1.23 ;
      POLYGON 8.02 1.11 4.82 1.11 4.82 1.43 4.34 1.43 4.34 1.55 4.46 1.55 4.46 1.67 4.22 1.67 4.22 1.43 2.87 1.43 2.87 1.19 2.99 1.19 2.99 1.31 4.7 1.31 4.7 0.71 4.72 0.71 4.72 0.59 4.84 0.59 4.84 0.83 4.82 0.83 4.82 0.99 8.02 0.99 ;
      POLYGON 4.56 1.19 4.02 1.19 4.02 1.07 4.44 1.07 4.44 0.95 4.06 0.95 4.06 0.48 3.45 0.48 3.45 0.83 2.43 0.83 2.43 1.79 2.55 1.79 2.55 1.91 2.31 1.91 2.31 0.61 2.33 0.61 2.33 0.49 2.45 0.49 2.45 0.71 3.33 0.71 3.33 0.36 4.18 0.36 4.18 0.83 4.56 0.83 ;
      POLYGON 3.59 2.11 3.35 2.11 3.35 1.91 2.95 1.91 2.95 2.15 2.71 2.15 2.71 2.25 2.47 2.25 2.47 2.15 2.07 2.15 2.07 2.09 1.54 2.09 1.54 1.86 1.4 1.86 1.4 1.5 1.555 1.5 1.555 0.86 1.46 0.86 1.46 0.74 1.7 0.74 1.7 0.86 1.675 0.86 1.675 1.62 1.52 1.62 1.52 1.74 1.66 1.74 1.66 1.97 2.07 1.97 2.07 0.85 2.19 0.85 2.19 2.03 2.83 2.03 2.83 1.79 3.47 1.79 3.47 1.99 3.59 1.99 ;
      POLYGON 2.03 0.73 1.95 0.73 1.95 1.85 1.83 1.85 1.83 0.62 1.21 0.62 1.21 0.68 0.68 0.68 0.68 0.92 0.53 0.92 0.53 1.575 0.46 1.575 0.46 1.695 0.34 1.695 0.34 1.455 0.41 1.455 0.41 0.8 0.56 0.8 0.56 0.56 1.09 0.56 1.09 0.5 1.91 0.5 1.91 0.49 2.03 0.49 ;
  END
END TLATNTSCAX20

MACRO AOI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21XL 0 0 ;
  SIZE 1.74 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.98 1.38 1.435 ;
        RECT 1.245 0.98 1.365 1.46 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 0.7 0.945 1.02 ;
        RECT 0.65 0.7 0.945 0.92 ;
        RECT 0.65 0.595 0.8 0.92 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.92 0.475 1.045 ;
        RECT 0.07 0.885 0.22 1.15 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.5 0.885 1.67 1.145 ;
        RECT 1.5 0.74 1.62 1.675 ;
        RECT 1.485 1.555 1.605 1.795 ;
        RECT 1.065 0.74 1.62 0.86 ;
        RECT 1.065 0.44 1.185 0.86 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.74 0.18 ;
        RECT 1.425 0.5 1.665 0.62 ;
        RECT 1.425 -0.18 1.545 0.62 ;
        RECT 0.345 -0.18 0.465 0.68 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.74 2.79 ;
        RECT 0.615 2.1 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.185 1.82 1.065 1.82 1.065 1.7 0.075 1.7 0.075 1.58 1.185 1.58 ;
  END
END AOI21XL

MACRO NAND2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX2 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.205 1.265 1.395 ;
        RECT 0.885 1.18 1.145 1.395 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 1.24 2.135 1.48 ;
        RECT 1.84 1.36 2.135 1.48 ;
        RECT 1.81 1.465 1.96 1.725 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.395 1.515 1.515 2.21 ;
        RECT 0.195 1.515 1.515 1.635 ;
        RECT 1.115 0.65 1.355 0.77 ;
        RECT 0.195 0.7 1.235 0.82 ;
        RECT 0.555 1.515 0.675 2.21 ;
        RECT 0.195 0.7 0.315 1.635 ;
        RECT 0.07 0.885 0.315 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.815 -0.18 1.935 0.64 ;
        RECT 0.475 0.46 0.715 0.58 ;
        RECT 0.475 -0.18 0.595 0.58 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.815 1.845 1.935 2.79 ;
        RECT 0.975 1.755 1.095 2.79 ;
        RECT 0.135 1.755 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.415 1.8 2.295 1.8 2.295 1.06 1.835 1.06 1.835 1.11 1.595 1.11 1.595 1.06 0.765 1.06 0.765 1.11 0.435 1.11 0.435 0.99 0.645 0.99 0.645 0.94 2.295 0.94 2.295 0.59 2.415 0.59 ;
  END
END NAND2BX2

MACRO NOR4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX4 0 0 ;
  SIZE 8.99 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.465 ;
        RECT 0.375 1.01 0.495 1.495 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 1.01 0.835 1.38 ;
        RECT 0.65 1.07 0.8 1.435 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.29 1.025 5.44 1.48 ;
        RECT 5.32 1 5.44 1.48 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.74 1.175 7.055 1.35 ;
        RECT 6.935 1.11 7.055 1.35 ;
        RECT 6.74 1.175 6.89 1.435 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.5168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.055 1.19 8.175 2.01 ;
        RECT 7.205 1.19 8.175 1.31 ;
        RECT 1.985 0.76 7.985 0.88 ;
        RECT 7.865 0.59 7.985 0.88 ;
        RECT 7.215 1.175 7.47 1.435 ;
        RECT 7.215 1.175 7.335 2.01 ;
        RECT 7.205 0.71 7.325 1.43 ;
        RECT 7.025 0.71 7.325 0.88 ;
        RECT 7.025 0.59 7.145 0.88 ;
        RECT 6.185 0.59 6.305 0.88 ;
        RECT 5.345 0.59 5.465 0.88 ;
        RECT 4.505 0.59 4.625 0.88 ;
        RECT 3.665 0.59 3.785 0.88 ;
        RECT 2.825 0.59 2.945 0.88 ;
        RECT 1.985 0.59 2.105 0.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.99 0.18 ;
        RECT 8.285 -0.18 8.405 0.64 ;
        RECT 7.445 -0.18 7.565 0.64 ;
        RECT 6.605 -0.18 6.725 0.64 ;
        RECT 5.765 -0.18 5.885 0.64 ;
        RECT 4.925 -0.18 5.045 0.64 ;
        RECT 4.085 -0.18 4.205 0.64 ;
        RECT 3.245 -0.18 3.365 0.64 ;
        RECT 2.405 -0.18 2.525 0.64 ;
        RECT 1.565 -0.18 1.685 0.64 ;
        RECT 0.555 -0.18 0.675 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.99 2.79 ;
        RECT 2.625 1.56 2.745 2.79 ;
        RECT 1.785 1.72 1.905 2.79 ;
        RECT 0.555 1.615 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.595 2.13 8.55 2.13 8.55 2.25 5.115 2.25 5.115 1.84 5.235 1.84 5.235 2.13 5.955 2.13 5.955 1.84 6.075 1.84 6.075 2.13 6.795 2.13 6.795 1.555 6.915 1.555 6.915 2.13 7.635 2.13 7.635 1.43 7.755 1.43 7.755 2.13 8.43 2.13 8.43 2.01 8.475 2.01 8.475 1.43 8.595 1.43 ;
      POLYGON 6.495 2.01 6.375 2.01 6.375 1.72 5.655 1.72 5.655 2.01 5.535 2.01 5.535 1.72 4.425 1.72 4.425 2.01 4.305 2.01 4.305 1.72 3.585 1.72 3.585 2.01 3.465 2.01 3.465 1.56 3.585 1.56 3.585 1.6 4.305 1.6 4.305 1.56 4.425 1.56 4.425 1.6 6.375 1.6 6.375 1.43 6.495 1.43 ;
      POLYGON 4.845 2.21 4.8 2.21 4.8 2.25 3.09 2.25 3.09 2.21 3.045 2.21 3.045 1.44 2.37 1.44 2.37 1.6 2.325 1.6 2.325 2.21 2.205 2.21 2.205 1.6 1.485 1.6 1.485 2.21 1.365 2.21 1.365 1.48 2.25 1.48 2.25 1.32 3.165 1.32 3.165 2.09 3.21 2.09 3.21 2.13 3.885 2.13 3.885 1.84 4.005 1.84 4.005 2.13 4.68 2.13 4.68 2.09 4.725 2.09 4.725 1.84 4.845 1.84 ;
      POLYGON 3.585 1.12 1.745 1.12 1.745 0.88 1.325 0.88 1.325 0.48 0.915 0.48 0.915 0.89 0.24 0.89 0.24 1.585 0.255 1.585 0.255 2.21 0.135 2.21 0.135 1.705 0.12 1.705 0.12 0.72 0.135 0.72 0.135 0.6 0.255 0.6 0.255 0.77 0.795 0.77 0.795 0.36 1.445 0.36 1.445 0.76 1.865 0.76 1.865 1 3.585 1 ;
      POLYGON 1.905 1.36 1.155 1.36 1.155 1.48 1.095 1.48 1.095 2.21 0.975 2.21 0.975 1.36 1.035 1.36 1.035 0.6 1.155 0.6 1.155 1.24 1.905 1.24 ;
  END
END NOR4BBX4

MACRO SDFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRXL 0 0 ;
  SIZE 12.76 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1.505 2.175 1.73 ;
        RECT 1.755 1.42 2.015 1.67 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.925 2.11 7.805 2.23 ;
        RECT 6.925 1.8 7.045 2.23 ;
        RECT 5.295 1.8 7.045 1.92 ;
        RECT 5.295 1.44 5.415 1.92 ;
        RECT 3.565 1.44 5.415 1.56 ;
        RECT 3.565 1.23 3.755 1.56 ;
        RECT 3.445 1.26 3.755 1.38 ;
        RECT 3.495 1.23 3.755 1.38 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.055 1.52 10.585 1.64 ;
        RECT 10.055 1.52 10.475 1.67 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.805 1.24 10.925 1.48 ;
        RECT 10.455 1.24 10.925 1.38 ;
        RECT 10.455 1.23 10.715 1.38 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.845 1.22 12.18 1.43 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 0.94 12.455 1.09 ;
        RECT 12.3 0.87 12.42 1.11 ;
        RECT 11.285 0.98 12.42 1.1 ;
        RECT 11.605 0.85 11.725 1.1 ;
        RECT 11.285 0.98 11.405 1.67 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.15 1.34 0.27 1.58 ;
        RECT 0.135 0.68 0.255 0.96 ;
        RECT 0.13 0.84 0.25 1.46 ;
        RECT 0.07 0.885 0.25 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 1.585 1.535 2.09 ;
        RECT 1.415 0.68 1.535 0.96 ;
        RECT 1.23 1.465 1.495 1.725 ;
        RECT 1.375 0.84 1.495 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 12.76 0.18 ;
        RECT 12.085 -0.18 12.205 0.75 ;
        RECT 10.685 0.5 10.925 0.62 ;
        RECT 10.805 -0.18 10.925 0.62 ;
        RECT 9.695 -0.18 9.935 0.32 ;
        RECT 7.825 -0.18 7.945 0.86 ;
        RECT 3.125 -0.18 3.365 0.32 ;
        RECT 1.835 -0.18 1.955 0.92 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 12.76 2.79 ;
        RECT 12.085 1.97 12.205 2.79 ;
        RECT 10.745 2.03 10.985 2.15 ;
        RECT 10.745 2.03 10.865 2.79 ;
        RECT 9.875 2.03 10.115 2.15 ;
        RECT 9.875 2.03 9.995 2.79 ;
        RECT 7.945 2.23 8.065 2.79 ;
        RECT 6.225 2.29 6.465 2.79 ;
        RECT 4.445 2.16 4.685 2.28 ;
        RECT 4.445 2.16 4.565 2.79 ;
        RECT 3.185 2.17 3.305 2.79 ;
        RECT 1.835 1.97 1.955 2.79 ;
        RECT 0.57 1.46 0.69 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 12.695 1.79 12.625 1.79 12.625 2.09 12.505 2.09 12.505 1.67 11.605 1.67 11.605 1.43 11.725 1.43 11.725 1.55 12.575 1.55 12.575 0.69 12.445 0.69 12.445 0.57 12.695 0.57 ;
      POLYGON 11.625 0.69 11.43 0.69 11.43 0.86 11.165 0.86 11.165 1.79 11.565 1.79 11.565 2.09 11.445 2.09 11.445 1.91 11.045 1.91 11.045 0.86 10.445 0.86 10.445 0.56 9.005 0.56 9.005 0.74 9.065 0.74 9.065 1.58 9.185 1.58 9.185 1.82 9.065 1.82 9.065 1.7 8.945 1.7 8.945 0.86 8.885 0.86 8.885 0.44 10.565 0.44 10.565 0.74 11.31 0.74 11.31 0.57 11.625 0.57 ;
      POLYGON 10.505 2.09 10.385 2.09 10.385 1.91 9.67 1.91 9.67 2.06 8.685 2.06 8.685 2.2 8.445 2.2 8.445 2.06 7.96 2.06 7.96 1.99 7.165 1.99 7.165 1.6 6.735 1.6 6.735 1.41 6.615 1.41 6.615 1.29 6.855 1.29 6.855 1.48 7.285 1.48 7.285 1.87 8.08 1.87 8.08 1.94 9.55 1.94 9.55 1.79 9.815 1.79 9.815 1.11 9.665 1.11 9.665 1.2 9.545 1.2 9.545 0.96 9.665 0.96 9.665 0.99 10.085 0.99 10.085 0.68 10.325 0.68 10.325 0.8 10.205 0.8 10.205 1.11 9.935 1.11 9.935 1.79 10.505 1.79 ;
      POLYGON 9.635 1.67 9.305 1.67 9.305 1.4 9.185 1.4 9.185 1.16 9.215 1.16 9.215 0.68 9.455 0.68 9.455 0.8 9.335 0.8 9.335 1.28 9.425 1.28 9.425 1.55 9.635 1.55 ;
      POLYGON 8.825 1.76 8.585 1.76 8.585 1.12 7.265 1.12 7.265 1 8.465 1 8.465 0.62 8.585 0.62 8.585 1 8.705 1 8.705 1.64 8.825 1.64 ;
      POLYGON 8.145 1.36 7.525 1.36 7.525 1.63 7.645 1.63 7.645 1.75 7.405 1.75 7.405 1.36 6.985 1.36 6.985 1.04 6.495 1.04 6.495 1.68 5.955 1.68 5.955 1.56 6.375 1.56 6.375 1.04 6.055 1.04 6.055 0.66 6.175 0.66 6.175 0.92 6.985 0.92 6.985 0.62 7.105 0.62 7.105 1.24 8.145 1.24 ;
      POLYGON 7.525 0.86 7.405 0.86 7.405 0.62 7.225 0.62 7.225 0.5 6.745 0.5 6.745 0.8 6.505 0.8 6.505 0.68 6.625 0.68 6.625 0.38 7.345 0.38 7.345 0.5 7.525 0.5 ;
      POLYGON 6.805 2.17 6.55 2.17 6.55 2.16 4.96 2.16 4.96 2.04 4.285 2.04 4.285 2.25 4.165 2.25 4.165 2.04 3.17 2.04 3.17 2.05 2.375 2.05 2.375 2.09 2.255 2.09 2.255 1.85 2.315 1.85 2.315 0.68 2.435 0.68 2.435 1.93 3.05 1.93 3.05 1.92 5.08 1.92 5.08 2.04 6.67 2.04 6.67 2.05 6.805 2.05 ;
      POLYGON 6.255 1.36 5.815 1.36 5.815 0.52 5.375 0.52 5.375 0.4 5.935 0.4 5.935 1.24 6.255 1.24 ;
      POLYGON 5.775 1.68 5.535 1.68 5.535 1.56 5.575 1.56 5.575 1.32 4.225 1.32 4.225 1.11 3.325 1.11 3.325 1.18 2.905 1.18 2.905 1.06 3.205 1.06 3.205 0.99 4.345 0.99 4.345 1.2 5.575 1.2 5.575 0.66 5.695 0.66 5.695 1.56 5.775 1.56 ;
      POLYGON 5.275 0.9 5.185 0.9 5.185 1.08 4.465 1.08 4.465 0.84 4.285 0.84 4.285 0.72 4.585 0.72 4.585 0.96 5.065 0.96 5.065 0.78 5.155 0.78 5.155 0.66 5.275 0.66 ;
      RECT 3.605 1.68 5.175 1.8 ;
      POLYGON 4.945 0.84 4.705 0.84 4.705 0.6 4.165 0.6 4.165 0.76 3.845 0.76 3.845 0.84 3.605 0.84 3.605 0.72 3.725 0.72 3.725 0.64 4.045 0.64 4.045 0.48 4.825 0.48 4.825 0.72 4.945 0.72 ;
      POLYGON 3.925 0.52 3.605 0.52 3.605 0.56 2.825 0.56 2.825 0.9 2.785 0.9 2.785 1.57 2.825 1.57 2.825 1.81 2.705 1.81 2.705 1.69 2.665 1.69 2.665 0.78 2.705 0.78 2.705 0.56 2.195 0.56 2.195 1.2 1.615 1.2 1.615 1.08 2.075 1.08 2.075 0.44 3.485 0.44 3.485 0.4 3.925 0.4 ;
      POLYGON 1.145 1.08 1.11 1.08 1.11 1.58 0.99 1.58 0.99 1.2 0.37 1.2 0.37 1.08 0.99 1.08 0.99 0.96 1.025 0.96 1.025 0.68 1.145 0.68 ;
  END
END SDFFSRXL

MACRO OR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1 0.51 1.455 ;
        RECT 0.375 1 0.495 1.485 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1 0.815 1.46 ;
        RECT 0.65 1 0.815 1.435 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.94 1.435 1.21 ;
        RECT 1.175 0.94 1.415 1.22 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 0.885 1.96 1.145 ;
        RECT 1.815 0.59 1.935 1.145 ;
        RECT 1.795 1.145 1.93 1.265 ;
        RECT 1.795 1.145 1.915 1.99 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.335 0.46 1.575 0.58 ;
        RECT 1.335 -0.18 1.455 0.58 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.375 1.34 1.495 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.675 1.17 1.555 1.17 1.555 0.82 1.055 0.82 1.055 1.725 0.155 1.725 0.155 1.605 0.935 1.605 0.935 0.88 0.135 0.88 0.135 0.4 0.255 0.4 0.255 0.76 0.935 0.76 0.935 0.7 0.975 0.7 0.975 0.4 1.095 0.4 1.095 0.7 1.675 0.7 ;
  END
END OR3X1

MACRO EDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRXL 0 0 ;
  SIZE 11.89 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.935 1.02 2.055 1.305 ;
        RECT 1.81 0.885 1.96 1.185 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.61 1.465 7.76 1.725 ;
        RECT 7.61 1.33 7.73 1.725 ;
        RECT 7.375 1.33 7.73 1.45 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.165 1.52 10.425 1.67 ;
        RECT 10.165 1.29 10.385 1.67 ;
        RECT 9.505 1.29 10.385 1.41 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.09 1.175 11.29 1.45 ;
        RECT 11.055 1.04 11.225 1.3 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 0.68 1.485 1.58 ;
        RECT 1.23 1.175 1.485 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.89 0.18 ;
        RECT 10.965 -0.18 11.085 0.92 ;
        RECT 9.345 0.57 9.585 0.69 ;
        RECT 9.345 -0.18 9.465 0.69 ;
        RECT 8.815 0.57 9.055 0.69 ;
        RECT 8.815 -0.18 8.935 0.69 ;
        RECT 7.695 0.6 7.935 0.72 ;
        RECT 7.815 -0.18 7.935 0.72 ;
        RECT 6.285 -0.18 6.525 0.32 ;
        RECT 4.685 0.65 4.925 0.77 ;
        RECT 4.685 -0.18 4.805 0.77 ;
        RECT 3.085 -0.18 3.205 0.38 ;
        RECT 1.845 -0.18 1.965 0.4 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.89 2.79 ;
        RECT 11.025 1.96 11.145 2.79 ;
        RECT 7.615 2.23 7.735 2.79 ;
        RECT 6.205 2.17 6.445 2.29 ;
        RECT 6.205 2.17 6.325 2.79 ;
        RECT 4.565 2.17 4.805 2.29 ;
        RECT 4.565 2.17 4.685 2.79 ;
        RECT 2.925 1.89 3.205 2.01 ;
        RECT 3.085 1.75 3.205 2.01 ;
        RECT 2.925 1.89 3.045 2.79 ;
        RECT 1.845 1.98 1.965 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.625 1.84 10.88 1.84 10.88 1.91 10.615 1.91 10.615 2.23 9.845 2.23 9.845 2.11 10.495 2.11 10.495 1.79 10.76 1.79 10.76 1.72 11.505 1.72 11.505 0.92 11.385 0.92 11.385 0.68 11.505 0.68 11.505 0.8 11.625 0.8 ;
      POLYGON 10.665 1.6 10.545 1.6 10.545 1.17 8.595 1.17 8.595 1.05 10.545 1.05 10.545 0.68 10.665 0.68 ;
      POLYGON 10.225 1.91 9.925 1.91 9.925 1.67 9.325 1.67 9.325 1.85 9.205 1.85 9.205 1.41 8.355 1.41 8.355 0.96 7.455 0.96 7.455 0.48 6.765 0.48 6.765 0.56 6.045 0.56 6.045 0.52 5.925 0.52 5.925 0.4 6.165 0.4 6.165 0.44 6.645 0.44 6.645 0.36 7.575 0.36 7.575 0.84 8.175 0.84 8.175 0.54 8.295 0.54 8.295 0.66 8.475 0.66 8.475 0.81 9.78 0.81 9.78 0.63 10.045 0.63 10.045 0.51 10.165 0.51 10.165 0.75 9.9 0.75 9.9 0.93 8.475 0.93 8.475 1.29 9.325 1.29 9.325 1.55 10.045 1.55 10.045 1.79 10.225 1.79 ;
      POLYGON 9.805 1.91 9.685 1.91 9.685 2.09 8.455 2.09 8.455 1.89 8.335 1.89 8.335 1.77 8.575 1.77 8.575 1.97 9.565 1.97 9.565 1.79 9.805 1.79 ;
      POLYGON 8.935 1.83 8.815 1.83 8.815 1.65 8.095 1.65 8.095 1.83 7.975 1.83 7.975 1.53 8.935 1.53 ;
      POLYGON 8.295 2.21 8.055 2.21 8.055 2.07 6.73 2.07 6.73 2.05 6.055 2.05 6.055 2.11 4.925 2.11 4.925 2.05 4.25 2.05 4.25 2.11 3.445 2.11 3.445 2.25 3.165 2.25 3.165 2.13 3.325 2.13 3.325 1.63 2.915 1.63 2.915 1.77 2.785 1.77 2.785 1.87 2.665 1.87 2.665 1.86 1.685 1.86 1.685 1.96 1.445 1.96 1.445 1.84 1.565 1.84 1.565 1.74 2.625 1.74 2.625 0.9 2.605 0.9 2.605 0.66 2.725 0.66 2.725 0.78 2.745 0.78 2.745 1.51 3.445 1.51 3.445 1.99 4.13 1.99 4.13 1.93 5.045 1.93 5.045 1.99 5.935 1.99 5.935 1.93 6.85 1.93 6.85 1.95 8.175 1.95 8.175 2.09 8.295 2.09 ;
      POLYGON 7.975 1.2 7.255 1.2 7.255 1.83 7.135 1.83 7.135 0.72 7.095 0.72 7.095 0.6 7.335 0.6 7.335 0.72 7.255 0.72 7.255 1.08 7.975 1.08 ;
      POLYGON 6.945 0.84 6.885 0.84 6.885 1.69 6.925 1.69 6.925 1.81 6.685 1.81 6.685 1.69 6.765 1.69 6.765 1.48 5.645 1.48 5.645 1.36 6.765 1.36 6.765 0.84 6.705 0.84 6.705 0.72 6.945 0.72 ;
      POLYGON 6.645 1.16 5.685 1.16 5.685 0.54 5.285 0.54 5.285 1.53 5.165 1.53 5.165 1.01 4.445 1.01 4.445 0.54 4.085 0.54 4.085 1.55 3.965 1.55 3.965 0.54 3.445 0.54 3.445 0.62 2.845 0.62 2.845 0.54 2.435 0.54 2.435 0.68 2.335 0.68 2.335 0.8 2.395 0.8 2.395 1.58 2.275 1.58 2.275 0.92 2.215 0.92 2.215 0.56 2.315 0.56 2.315 0.42 2.965 0.42 2.965 0.5 3.325 0.5 3.325 0.42 3.445 0.42 3.445 0.38 3.685 0.38 3.685 0.42 4.565 0.42 4.565 0.89 5.165 0.89 5.165 0.42 5.805 0.42 5.805 1.04 6.645 1.04 ;
      POLYGON 5.565 1.24 5.525 1.24 5.525 1.87 5.405 1.87 5.405 1.77 4.925 1.77 4.925 1.49 4.445 1.49 4.445 1.37 5.045 1.37 5.045 1.65 5.405 1.65 5.405 1.12 5.445 1.12 5.445 0.66 5.565 0.66 ;
      POLYGON 5.025 1.25 4.325 1.25 4.325 1.81 4.085 1.81 4.085 1.69 4.205 1.69 4.205 0.66 4.325 0.66 4.325 1.13 5.025 1.13 ;
      POLYGON 3.845 1.87 3.725 1.87 3.725 1.39 2.865 1.39 2.865 1.27 3.725 1.27 3.725 0.84 3.605 0.84 3.605 0.72 3.845 0.72 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END EDFFTRXL

MACRO BUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX6 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 1.39 2.01 2.21 ;
        RECT 0.15 0.91 2.01 1.03 ;
        RECT 1.89 0.4 2.01 1.03 ;
        RECT 0.21 1.39 2.01 1.51 ;
        RECT 1.05 1.39 1.17 2.21 ;
        RECT 0.99 0.4 1.11 1.03 ;
        RECT 0.36 1.175 0.51 1.51 ;
        RECT 0.36 0.91 0.48 1.51 ;
        RECT 0.21 1.39 0.33 2.21 ;
        RECT 0.15 0.4 0.27 1.03 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.825 3.12 1.285 ;
        RECT 2.97 0.825 3.09 1.31 ;
    END
  END A
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 3.15 1.43 3.27 2.79 ;
        RECT 2.31 1.43 2.43 2.79 ;
        RECT 1.47 1.63 1.59 2.79 ;
        RECT 0.63 1.63 0.75 2.79 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 3.15 -0.18 3.27 0.705 ;
        RECT 2.31 -0.18 2.43 0.895 ;
        RECT 1.41 -0.18 1.53 0.79 ;
        RECT 0.57 -0.18 0.69 0.79 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.85 2.08 2.73 2.08 2.73 1.27 0.77 1.27 0.77 1.15 2.73 1.15 2.73 0.655 2.85 0.655 ;
  END
END BUFX6

MACRO NOR3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BXL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1 0.51 1.5 ;
        RECT 0.36 1 0.51 1.47 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.935 1.4 ;
        RECT 0.815 1.16 0.935 1.4 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.465 1.15 1.725 1.38 ;
        RECT 1.475 1.09 1.595 1.5 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2448 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 0.46 1.155 0.58 ;
        RECT 0.12 0.76 1.035 0.88 ;
        RECT 0.915 0.46 1.035 0.88 ;
        RECT 0.335 1.62 0.455 1.86 ;
        RECT 0.12 1.62 0.455 1.74 ;
        RECT 0.135 0.4 0.255 0.88 ;
        RECT 0.12 0.76 0.24 1.74 ;
        RECT 0.07 0.885 0.24 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.395 -0.18 1.515 0.64 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.295 1.62 1.415 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.965 1.62 1.835 1.62 1.835 1.74 1.715 1.74 1.715 1.5 1.845 1.5 1.845 0.97 1.345 0.97 1.345 1.06 1.225 1.06 1.225 0.82 1.345 0.82 1.345 0.85 1.845 0.85 1.845 0.64 1.815 0.64 1.815 0.4 1.935 0.4 1.935 0.52 1.965 0.52 ;
  END
END NOR3BXL

MACRO MXI3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X1 0 0 ;
  SIZE 6.09 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.52 1.455 1.64 ;
        RECT 1.335 1.36 1.455 1.64 ;
        RECT 0.305 1.52 0.565 1.67 ;
        RECT 0.355 1.34 0.475 1.67 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.21 1.035 1.365 ;
        RECT 0.595 1.21 0.855 1.4 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.5 2.595 1.67 ;
        RECT 2.255 1.34 2.375 1.62 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.455 1.4 4.475 1.52 ;
        RECT 3.455 1.23 3.755 1.52 ;
        RECT 3.455 1.16 3.695 1.52 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 0.9 5.205 1.115 ;
        RECT 4.965 0.9 5.085 1.28 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.665 0.68 5.785 1.99 ;
        RECT 5.58 0.885 5.785 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.09 0.18 ;
        RECT 5.245 -0.18 5.365 0.78 ;
        RECT 3.955 0.68 4.195 0.8 ;
        RECT 3.955 -0.18 4.075 0.8 ;
        RECT 2.275 -0.18 2.395 0.86 ;
        RECT 0.655 0.68 0.895 0.8 ;
        RECT 0.655 -0.18 0.775 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.09 2.79 ;
        RECT 5.125 1.88 5.365 2 ;
        RECT 5.125 1.88 5.245 2.79 ;
        RECT 3.695 2.22 3.935 2.79 ;
        RECT 2.335 1.8 2.455 2.79 ;
        RECT 0.795 1.8 0.915 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.46 1.52 5.215 1.52 5.215 1.76 4.95 1.76 4.95 2.1 2.975 2.1 2.975 1.86 2.855 1.86 2.855 0.68 3.095 0.68 3.095 0.8 2.975 0.8 2.975 1.74 3.095 1.74 3.095 1.98 4.83 1.98 4.83 1.64 5.095 1.64 5.095 1.4 5.34 1.4 5.34 1.02 5.46 1.02 ;
      POLYGON 4.945 0.78 4.795 0.78 4.795 1.28 4.765 1.28 4.765 1.4 4.885 1.4 4.885 1.52 4.645 1.52 4.645 1.28 3.875 1.28 3.875 1.16 4.675 1.16 4.675 0.66 4.825 0.66 4.825 0.54 4.945 0.54 ;
      POLYGON 4.555 1.04 3.64 1.04 3.64 0.56 3.335 0.56 3.335 1.64 4.295 1.64 4.295 1.74 4.415 1.74 4.415 1.86 4.175 1.86 4.175 1.76 3.215 1.76 3.215 1.54 3.095 1.54 3.095 1.42 3.215 1.42 3.215 0.56 3.1 0.56 3.1 0.48 2.715 0.48 2.715 0.36 3.22 0.36 3.22 0.44 3.76 0.44 3.76 0.92 4.435 0.92 4.435 0.62 4.555 0.62 ;
      POLYGON 2.555 1.22 2.135 1.22 2.135 1.82 1.795 1.82 1.795 1.88 1.555 1.88 1.555 1.76 1.675 1.76 1.675 1.7 2.015 1.7 2.015 1.22 1.815 1.22 1.815 0.8 1.295 0.8 1.295 0.68 1.935 0.68 1.935 1.1 2.435 1.1 2.435 0.98 2.555 0.98 ;
      POLYGON 1.895 1.58 1.775 1.58 1.775 1.46 1.575 1.46 1.575 1.12 1.155 1.12 1.155 1.09 0.185 1.09 0.185 1.79 0.495 1.79 0.495 2.03 0.375 2.03 0.375 1.91 0.065 1.91 0.065 0.74 0.295 0.74 0.295 0.62 0.415 0.62 0.415 0.97 1.695 0.97 1.695 1.34 1.895 1.34 ;
  END
END MXI3X1

MACRO NAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.99 3.315 1.11 ;
        RECT 0.595 0.94 0.855 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.335 1.23 2.595 1.38 ;
        RECT 1.175 1.23 2.595 1.35 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1072 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.5 3.555 1.62 ;
        RECT 3.435 0.7 3.555 1.62 ;
        RECT 3.205 1.23 3.555 1.38 ;
        RECT 1.335 0.7 3.555 0.82 ;
        RECT 3.075 1.5 3.195 2.21 ;
        RECT 2.495 0.65 2.735 0.82 ;
        RECT 2.235 1.5 2.355 2.21 ;
        RECT 1.395 1.5 1.515 2.21 ;
        RECT 1.215 0.65 1.455 0.77 ;
        RECT 0.555 1.5 0.675 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.135 0.46 3.375 0.58 ;
        RECT 3.135 -0.18 3.255 0.58 ;
        RECT 1.855 0.46 2.095 0.58 ;
        RECT 1.855 -0.18 1.975 0.58 ;
        RECT 0.635 -0.18 0.755 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.56 0.255 2.79 ;
    END
  END VDD
END NAND2X4

MACRO AOI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X1 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.78 0.51 1.215 ;
        RECT 0.38 0.78 0.5 1.32 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.135 1.025 2.54 1.145 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.135 1.025 2.255 1.265 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.04 0.82 1.16 1.17 ;
        RECT 0.94 0.595 1.09 0.945 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.94 2.015 1.095 ;
        RECT 1.52 0.985 1.875 1.11 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.845 0.82 1.27 ;
        RECT 0.65 0.56 0.8 0.965 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3778 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.26 1.935 2.01 ;
        RECT 1.28 1.26 1.935 1.38 ;
        RECT 1.28 1.23 1.725 1.38 ;
        RECT 1.32 0.61 1.44 0.865 ;
        RECT 1.28 0.745 1.4 1.38 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 2.08 -0.18 2.2 0.66 ;
        RECT 0.22 -0.18 0.34 0.66 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.5 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.355 2.25 1.395 2.25 1.395 1.62 0.675 1.62 0.675 2.15 0.555 2.15 0.555 1.5 1.515 1.5 1.515 2.13 2.235 2.13 2.235 1.5 2.355 1.5 ;
  END
END AOI32X1

MACRO NAND4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX1 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.785 0.51 1.24 ;
        RECT 0.39 0.76 0.51 1.24 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.89 0.93 1.01 1.17 ;
        RECT 0.65 0.93 1.01 1.145 ;
        RECT 0.65 0.885 0.8 1.145 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.885 1.415 1.215 ;
        RECT 1.21 0.845 1.365 1.17 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 1 2.25 1.47 ;
        RECT 2.1 1 2.22 1.5 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5364 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.47 1.36 1.59 2.21 ;
        RECT 0.12 1.36 1.59 1.48 ;
        RECT 0.63 1.36 0.75 2.21 ;
        RECT 0.12 0.52 0.53 0.64 ;
        RECT 0.41 0.4 0.53 0.64 ;
        RECT 0.07 1.175 0.24 1.435 ;
        RECT 0.12 0.52 0.24 1.48 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.69 -0.18 1.81 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.89 1.62 2.01 2.79 ;
        RECT 1.05 1.6 1.17 2.79 ;
        RECT 0.21 1.6 0.33 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.49 1.8 2.37 1.8 2.37 0.88 1.98 0.88 1.98 1.11 1.63 1.11 1.63 0.99 1.86 0.99 1.86 0.76 2.17 0.76 2.17 0.59 2.29 0.59 2.29 0.71 2.49 0.71 ;
  END
END NAND4BX1

MACRO AO22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.885 0.82 1.32 ;
        RECT 0.7 0.86 0.82 1.32 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.98 1.09 1.16 1.33 ;
        RECT 0.94 1.175 1.145 1.435 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.03 0.51 1.5 ;
        RECT 0.36 1.03 0.48 1.53 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 1.96 1.81 ;
        RECT 1.52 1.465 1.96 1.585 ;
        RECT 1.52 1.41 1.8 1.585 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.4 2.825 1.52 ;
        RECT 2.39 0.885 2.54 1.145 ;
        RECT 2.39 0.885 2.51 1.52 ;
        RECT 2.16 0.885 2.54 1.025 ;
        RECT 2.16 0.67 2.28 1.025 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.68 0.73 1.92 0.85 ;
        RECT 1.68 -0.18 1.8 0.85 ;
        RECT 0.2 -0.18 0.32 0.91 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 2.205 1.98 2.325 2.79 ;
        RECT 0.555 1.89 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.04 1.31 1.92 1.31 1.92 1.29 1.4 1.29 1.4 1.705 1.515 1.705 1.515 2.01 1.395 2.01 1.395 1.825 1.28 1.825 1.28 0.97 1.06 0.97 1.06 0.85 0.94 0.85 0.94 0.73 1.18 0.73 1.18 0.85 1.4 0.85 1.4 1.17 1.92 1.17 1.92 1.07 2.04 1.07 ;
      POLYGON 1.995 2.07 1.875 2.07 1.875 2.25 0.975 2.25 0.975 1.77 0.315 1.77 0.315 1.95 0.075 1.95 0.075 1.83 0.195 1.83 0.195 1.65 1.095 1.65 1.095 2.13 1.755 2.13 1.755 1.95 1.995 1.95 ;
  END
END AO22XL

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.535 0.99 1.775 1.11 ;
        RECT 0.595 0.94 1.655 0.99 ;
        RECT 0.735 0.87 1.655 0.99 ;
        RECT 0.575 0.99 0.855 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 1.11 1.38 1.58 ;
        RECT 1.23 1.11 1.35 1.61 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.695 1.73 2.015 1.85 ;
        RECT 1.895 0.63 2.015 1.85 ;
        RECT 1.755 1.23 2.015 1.38 ;
        RECT 1.055 0.63 2.015 0.75 ;
        RECT 1.535 1.56 1.655 2.21 ;
        RECT 0.695 1.56 0.815 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.755 0.39 1.995 0.51 ;
        RECT 1.755 -0.18 1.875 0.51 ;
        RECT 0.475 -0.18 0.595 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.955 1.97 2.075 2.79 ;
        RECT 1.115 1.97 1.235 2.79 ;
        RECT 0.275 1.56 0.395 2.79 ;
    END
  END VDD
END NAND2X2

MACRO NOR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.06 1.8 1.22 ;
        RECT 1.52 1.1 1.67 1.435 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.28 1.05 1.4 1.475 ;
        RECT 1.23 1.175 1.38 1.585 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.05 1.09 1.505 ;
        RECT 0.96 1.05 1.08 1.535 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.13 0.615 1.3 ;
        RECT 0.295 1.18 0.565 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2544 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.92 0.81 2.04 1.585 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 0.7 0.81 2.04 0.93 ;
        RECT 1.79 1.465 1.96 1.705 ;
        RECT 1.54 0.45 1.66 0.93 ;
        RECT 0.7 0.45 0.82 0.93 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.96 -0.18 2.08 0.69 ;
        RECT 1.12 -0.18 1.24 0.69 ;
        RECT 0.28 -0.18 0.4 0.69 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 0.48 1.51 0.6 2.79 ;
    END
  END VDD
END NOR4XL

MACRO MX3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3XL 0 0 ;
  SIZE 4.93 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.71 1.25 0.83 1.555 ;
        RECT 0.65 1.435 0.8 1.75 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.785 2.54 1.18 ;
        RECT 2.38 1.06 2.5 1.47 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.72 0.785 2.84 1.27 ;
        RECT 2.68 0.77 2.83 1.23 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.8 1.01 4.04 1.13 ;
        RECT 3.84 1.01 3.99 1.435 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.13 1.465 4.28 1.725 ;
        RECT 4.14 1.435 4.26 1.725 ;
        RECT 3.56 1.555 4.28 1.675 ;
        RECT 3.56 1.25 3.68 1.675 ;
        RECT 3.48 1.11 3.6 1.37 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.17 1.85 0.41 1.97 ;
        RECT 0.29 0.61 0.41 1.97 ;
        RECT 0.07 0.885 0.41 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.93 0.18 ;
        RECT 3.98 -0.18 4.1 0.65 ;
        RECT 2.7 -0.18 2.82 0.65 ;
        RECT 0.71 -0.18 0.83 0.85 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.93 2.79 ;
        RECT 3.98 1.97 4.1 2.79 ;
        RECT 2.7 1.97 2.82 2.79 ;
        RECT 0.65 1.91 0.77 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.52 2.09 4.4 2.09 4.4 0.89 3.68 0.89 3.68 0.99 3.36 0.99 3.36 1.49 3.44 1.49 3.44 1.61 3.2 1.61 3.2 1.49 3.24 1.49 3.24 0.87 3.44 0.87 3.44 0.81 3.56 0.81 3.56 0.77 4.4 0.77 4.4 0.41 4.52 0.41 ;
      POLYGON 3.46 0.65 3.32 0.65 3.32 0.75 3.08 0.75 3.08 1.73 3.44 1.73 3.44 1.85 3.46 1.85 3.46 2.09 3.34 2.09 3.34 1.97 3.32 1.97 3.32 1.85 2.09 1.85 2.09 1.97 1.83 1.97 1.83 1.85 1.97 1.85 1.97 0.85 1.89 0.85 1.89 0.61 2.01 0.61 2.01 0.73 2.09 0.73 2.09 1.73 2.96 1.73 2.96 0.63 3.2 0.63 3.2 0.53 3.34 0.53 3.34 0.41 3.46 0.41 ;
      POLYGON 2.4 0.65 2.28 0.65 2.28 0.49 1.77 0.49 1.77 0.97 1.85 0.97 1.85 1.21 1.77 1.21 1.77 1.57 1.71 1.57 1.71 2.09 2.28 2.09 2.28 1.97 2.4 1.97 2.4 2.21 1.59 2.21 1.59 1.57 1.31 1.57 1.31 1.69 1.19 1.69 1.19 1.45 1.65 1.45 1.65 0.37 2.4 0.37 ;
      POLYGON 1.53 1.11 1.07 1.11 1.07 1.81 1.35 1.81 1.35 1.85 1.47 1.85 1.47 1.97 1.23 1.97 1.23 1.93 0.95 1.93 0.95 1.11 0.53 1.11 0.53 0.99 1.41 0.99 1.41 0.61 1.53 0.61 ;
  END
END MX3XL

MACRO CLKINVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX8 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.864 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.905 1.205 2.265 1.325 ;
        RECT 0.885 1.23 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.145 0.74 3.385 0.86 ;
        RECT 3.205 1.47 3.325 2.21 ;
        RECT 0.745 0.79 3.265 0.91 ;
        RECT 0.685 1.5 3.325 1.62 ;
        RECT 2.385 0.79 2.54 1.145 ;
        RECT 2.385 0.79 2.505 1.62 ;
        RECT 2.365 1.47 2.485 2.21 ;
        RECT 2.365 0.67 2.485 0.91 ;
        RECT 1.465 0.74 1.705 0.91 ;
        RECT 1.525 1.465 1.645 2.21 ;
        RECT 0.625 0.74 0.865 0.86 ;
        RECT 0.685 1.5 0.805 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.785 -0.18 2.905 0.67 ;
        RECT 1.945 -0.18 2.065 0.67 ;
        RECT 1.105 -0.18 1.225 0.67 ;
        RECT 0.265 -0.18 0.385 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.785 1.74 2.905 2.79 ;
        RECT 1.945 1.74 2.065 2.79 ;
        RECT 1.105 1.74 1.225 2.79 ;
        RECT 0.265 1.465 0.385 2.79 ;
    END
  END VDD
END CLKINVX8

MACRO OAI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1XL 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 0.885 1.67 1.355 ;
        RECT 1.55 0.855 1.67 1.355 ;
    END
  END A1N
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.16 1.53 ;
        RECT 1.04 1.17 1.16 1.53 ;
    END
  END A0N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.135 0.8 1.59 ;
        RECT 0.68 1.11 0.8 1.59 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1824 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.495 1.71 0.615 1.95 ;
        RECT 0.41 1.11 0.53 1.83 ;
        RECT 0.115 1.11 0.53 1.23 ;
        RECT 0.115 0.63 0.395 0.75 ;
        RECT 0.275 0.49 0.395 0.75 ;
        RECT 0.07 0.885 0.235 1.145 ;
        RECT 0.115 0.63 0.235 1.23 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 0.915 -0.18 1.035 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 2.23 1.895 2.79 ;
        RECT 0.975 2.23 1.095 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.675 0.735 1.4 0.735 1.4 1.475 1.455 1.475 1.455 1.83 1.335 1.83 1.335 1.595 1.28 1.595 1.28 0.99 0.355 0.99 0.355 0.87 1.28 0.87 1.28 0.615 1.555 0.615 1.555 0.49 1.675 0.49 ;
  END
END OAI2BB1XL

MACRO AOI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.66 0.82 1.105 ;
        RECT 0.65 0.72 0.8 1.145 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.115 0.885 1.235 1.245 ;
        RECT 0.94 0.885 1.235 1.24 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.815 1.125 1.935 1.52 ;
        RECT 1.465 1.155 1.935 1.38 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.29 0.885 0.53 1.09 ;
        RECT 0.36 0.885 0.51 1.28 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1992 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.055 1.175 2.25 1.435 ;
        RECT 2.055 0.885 2.175 1.685 ;
        RECT 1.375 0.885 2.175 1.005 ;
        RECT 1.375 0.525 1.495 1.005 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.795 -0.18 1.915 0.765 ;
        RECT 0.22 -0.18 0.34 0.765 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.095 2.085 1.215 2.79 ;
        RECT 0.135 2.085 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.695 1.745 1.575 1.745 1.575 1.625 0.555 1.625 0.555 1.505 1.695 1.505 ;
  END
END AOI31XL

MACRO DLY1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X1 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 1.175 0.8 1.435 ;
        RECT 0.395 1.18 0.8 1.42 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.735 0.67 2.855 2.21 ;
        RECT 2.68 0.885 2.855 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.315 -0.18 2.435 0.72 ;
        RECT 1.195 1.32 1.475 1.44 ;
        RECT 1.355 0.76 1.475 1.44 ;
        RECT 0.955 0.76 1.475 0.88 ;
        RECT 0.955 -0.18 1.075 0.88 ;
        RECT 0.555 -0.18 0.675 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.315 1.56 2.435 2.79 ;
        RECT 0.955 1 1.235 1.12 ;
        RECT 0.955 1 1.075 2.79 ;
        RECT 0.555 1.7 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.56 1.23 2.415 1.23 2.415 1.44 1.955 1.44 1.955 1.8 1.835 1.8 1.835 1.32 2.295 1.32 2.295 0.96 1.835 0.96 1.835 0.67 1.955 0.67 1.955 0.84 2.56 0.84 ;
      POLYGON 2.175 1.2 1.715 1.2 1.715 1.68 1.315 1.68 1.315 1.82 1.195 1.82 1.195 1.56 1.595 1.56 1.595 0.64 1.195 0.64 1.195 0.4 1.315 0.4 1.315 0.52 1.715 0.52 1.715 1.08 2.175 1.08 ;
      POLYGON 0.835 1 0.255 1 0.255 1.82 0.135 1.82 0.135 0.4 0.255 0.4 0.255 0.88 0.835 0.88 ;
  END
END DLY1X1

MACRO OAI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X4 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.055 1.23 4.755 1.35 ;
        RECT 4.055 1.23 4.335 1.38 ;
        RECT 4.055 1.195 4.175 1.435 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 1.175 3.41 1.435 ;
        RECT 3.235 0.99 3.38 1.23 ;
        RECT 0.615 0.99 3.38 1.11 ;
        RECT 1.775 0.99 2.015 1.16 ;
        RECT 0.495 1.02 0.735 1.14 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.195 1.28 2.655 1.4 ;
        RECT 1.175 1.23 1.435 1.38 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1072 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.775 0.7 5.015 0.82 ;
        RECT 3.815 0.81 4.895 0.93 ;
        RECT 4.635 1.555 4.755 2.21 ;
        RECT 1.355 1.555 4.755 1.675 ;
        RECT 3.815 0.7 4.175 0.93 ;
        RECT 3.795 1.555 3.99 2.015 ;
        RECT 3.815 0.7 3.935 2.015 ;
        RECT 3.795 1.555 3.915 2.21 ;
        RECT 2.635 1.555 2.755 2.21 ;
        RECT 1.355 1.555 1.475 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 3.095 0.51 3.335 0.63 ;
        RECT 3.095 -0.18 3.215 0.63 ;
        RECT 2.255 0.51 2.495 0.63 ;
        RECT 2.255 -0.18 2.375 0.63 ;
        RECT 1.415 0.51 1.655 0.63 ;
        RECT 1.415 -0.18 1.535 0.63 ;
        RECT 0.575 0.51 0.815 0.63 ;
        RECT 0.575 -0.18 0.695 0.63 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 5.055 1.56 5.175 2.79 ;
        RECT 4.215 1.795 4.335 2.79 ;
        RECT 3.375 1.795 3.495 2.79 ;
        RECT 1.995 1.795 2.115 2.79 ;
        RECT 0.415 1.56 0.535 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.375 0.7 5.255 0.7 5.255 0.58 4.535 0.58 4.535 0.69 4.415 0.69 4.415 0.58 3.695 0.58 3.695 0.87 0.215 0.87 0.215 0.63 0.335 0.63 0.335 0.75 1.055 0.75 1.055 0.63 1.175 0.63 1.175 0.75 1.895 0.75 1.895 0.63 2.015 0.63 2.015 0.75 2.735 0.75 2.735 0.63 2.855 0.63 2.855 0.75 3.575 0.75 3.575 0.46 4.415 0.46 4.415 0.45 4.535 0.45 4.535 0.46 5.375 0.46 ;
  END
END OAI21X4

MACRO SDFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX8 0 0 ;
  SIZE 13.92 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.775 0.665 2.895 0.96 ;
        RECT 2.655 0.84 2.775 2.085 ;
        RECT 0.255 1.025 2.775 1.145 ;
        RECT 1.935 0.665 2.055 1.145 ;
        RECT 1.815 0.905 1.935 2.085 ;
        RECT 1.095 0.665 1.215 1.145 ;
        RECT 0.975 0.905 1.095 2.08 ;
        RECT 0.255 0.885 0.51 1.145 ;
        RECT 0.255 0.665 0.375 1.265 ;
        RECT 0.135 1.145 0.255 2.08 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.402 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.41 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.9805 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.415 0.98 4.695 1.1 ;
        RECT 4.415 0.36 4.535 1.1 ;
        RECT 3.635 0.36 4.535 0.48 ;
        RECT 3.375 1 3.755 1.12 ;
        RECT 3.635 0.36 3.755 1.12 ;
        RECT 3.495 0.94 3.755 1.12 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.105 1.185 6.365 1.41 ;
        RECT 6.245 1.01 6.365 1.41 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.525 0.93 11.645 1.17 ;
        RECT 11.09 0.93 11.645 1.05 ;
        RECT 11.09 0.885 11.24 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.74 1.23 13.055 1.43 ;
        RECT 12.74 1.21 13.035 1.435 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.155 0.99 13.395 1.11 ;
        RECT 12.005 0.97 13.325 1.09 ;
        RECT 13.065 0.94 13.325 1.09 ;
        RECT 12.005 0.97 12.125 1.44 ;
    END
  END SE
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.92 0.18 ;
        RECT 13.065 -0.18 13.185 0.82 ;
        RECT 11.525 -0.18 11.645 0.64 ;
        RECT 8.585 0.43 8.825 0.55 ;
        RECT 8.705 -0.18 8.825 0.55 ;
        RECT 6.325 -0.18 6.565 0.41 ;
        RECT 4.755 -0.18 4.875 0.65 ;
        RECT 3.195 -0.18 3.315 0.65 ;
        RECT 2.355 -0.18 2.475 0.655 ;
        RECT 1.515 -0.18 1.635 0.655 ;
        RECT 0.675 -0.18 0.795 0.655 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.92 2.79 ;
        RECT 12.905 1.795 13.025 2.79 ;
        RECT 11.405 2.28 11.645 2.79 ;
        RECT 9.305 2.26 9.545 2.79 ;
        RECT 8.405 1.75 8.525 2.79 ;
        RECT 6.385 2.25 6.625 2.79 ;
        RECT 5.595 2.25 5.835 2.79 ;
        RECT 4.755 1.7 4.875 1.99 ;
        RECT 4.735 1.87 4.855 2.79 ;
        RECT 3.915 1.7 4.035 2.79 ;
        RECT 3.075 1.7 3.195 2.79 ;
        RECT 2.235 1.34 2.355 2.79 ;
        RECT 1.395 1.34 1.515 2.79 ;
        RECT 0.555 1.34 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.635 1.68 13.505 1.68 13.505 1.8 13.385 1.8 13.385 1.675 12.405 1.675 12.405 1.24 12.525 1.24 12.525 1.555 13.515 1.555 13.515 0.82 13.485 0.82 13.485 0.58 13.605 0.58 13.605 0.7 13.635 0.7 ;
      POLYGON 12.545 0.85 11.885 0.85 11.885 1.56 12.285 1.56 12.285 2.21 12.165 2.21 12.165 1.68 11.885 1.68 11.885 1.8 11.62 1.8 11.62 1.98 10.595 1.98 10.595 1.3 10.135 1.3 10.135 0.72 10.085 0.72 10.085 0.6 10.325 0.6 10.325 0.72 10.255 0.72 10.255 1.18 10.715 1.18 10.715 1.86 11.5 1.86 11.5 1.68 11.765 1.68 11.765 0.73 12.425 0.73 12.425 0.59 12.545 0.59 ;
      POLYGON 11.285 2.22 9.72 2.22 9.72 2.14 8.645 2.14 8.645 1.63 8.285 1.63 8.285 2.01 6.985 2.01 6.985 1.89 6.925 1.89 6.925 0.89 5.965 0.89 5.965 1.53 6.225 1.53 6.225 1.65 5.845 1.65 5.845 0.72 5.725 0.72 5.725 0.6 5.965 0.6 5.965 0.77 7.045 0.77 7.045 1.77 7.105 1.77 7.105 1.89 7.465 1.89 7.465 1.13 7.585 1.13 7.585 1.89 8.165 1.89 8.165 1.51 8.765 1.51 8.765 2.02 9.84 2.02 9.84 2.1 11.285 2.1 ;
      POLYGON 11.165 1.74 10.85 1.74 10.85 1.06 10.375 1.06 10.375 0.94 10.495 0.94 10.495 0.48 9.545 0.48 9.545 0.86 9.645 0.86 9.645 1.1 9.425 1.1 9.425 0.79 8.345 0.79 8.345 0.48 7.865 0.48 7.865 0.92 7.985 0.92 7.985 1.04 7.745 1.04 7.745 0.36 8.465 0.36 8.465 0.67 9.425 0.67 9.425 0.36 10.615 0.36 10.615 0.94 10.85 0.94 10.85 0.59 10.97 0.59 10.97 1.62 11.165 1.62 ;
      POLYGON 10.295 1.94 10.175 1.94 10.175 1.54 9.765 1.54 9.765 1.39 8.465 1.39 8.465 1.31 8.345 1.31 8.345 1.19 8.585 1.19 8.585 1.27 9.765 1.27 9.765 0.72 9.665 0.72 9.665 0.6 9.905 0.6 9.905 0.72 9.885 0.72 9.885 1.42 10.295 1.42 ;
      POLYGON 9.875 1.9 8.885 1.9 8.885 1.51 9.005 1.51 9.005 1.78 9.755 1.78 9.755 1.66 9.875 1.66 ;
      POLYGON 9.305 1.15 9.185 1.15 9.185 1.07 8.225 1.07 8.225 1.28 8.045 1.28 8.045 1.77 7.925 1.77 7.925 1.16 8.105 1.16 8.105 0.72 7.985 0.72 7.985 0.6 8.225 0.6 8.225 0.95 9.185 0.95 9.185 0.91 9.305 0.91 ;
      POLYGON 8.085 2.25 6.745 2.25 6.745 2.13 5.215 2.13 5.215 2.25 4.975 2.25 4.975 2.13 5.095 2.13 5.095 2.01 6.865 2.01 6.865 2.13 8.085 2.13 ;
      POLYGON 7.345 1.77 7.225 1.77 7.225 0.65 6.085 0.65 6.085 0.48 5.48 0.48 5.48 0.54 5.215 0.54 5.215 1.08 5.435 1.08 5.435 1.2 5.215 1.2 5.215 1.34 4.175 1.34 4.175 1 4.295 1 4.295 1.22 5.095 1.22 5.095 0.42 5.36 0.42 5.36 0.36 6.205 0.36 6.205 0.53 7.345 0.53 ;
      POLYGON 6.725 1.89 5.555 1.89 5.555 1.58 5.295 1.58 5.295 1.89 5.175 1.89 5.175 1.58 4.455 1.58 4.455 1.99 4.335 1.99 4.335 1.58 3.615 1.58 3.615 1.99 3.495 1.99 3.495 1.58 3.015 1.58 3.015 1.2 2.895 1.2 2.895 1.08 3.135 1.08 3.135 1.46 3.495 1.46 3.495 1.34 3.615 1.34 3.615 1.46 3.915 1.46 3.915 0.6 4.035 0.6 4.035 1.46 5.555 1.46 5.555 0.96 5.335 0.96 5.335 0.66 5.575 0.66 5.575 0.84 5.675 0.84 5.675 1.77 6.605 1.77 6.605 1.13 6.725 1.13 ;
  END
END SDFFRHQX8

MACRO NAND4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX2 0 0 ;
  SIZE 5.8 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.445 1.18 0.565 1.67 ;
        RECT 0.305 1.18 0.565 1.4 ;
    END
  END BN
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.52 1.145 1.705 ;
        RECT 0.885 1.33 1.005 1.705 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.095 1.03 4.28 1.435 ;
        RECT 4.095 1.015 4.215 1.435 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.815 1.075 4.935 1.38 ;
        RECT 4.71 0.88 4.86 1.195 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.9696 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.075 0.605 5.195 0.845 ;
        RECT 4.875 1.555 5.175 1.68 ;
        RECT 5.055 0.725 5.175 1.68 ;
        RECT 4.875 1.555 4.995 2.21 ;
        RECT 2.355 1.555 5.175 1.675 ;
        RECT 4.035 1.555 4.155 2.21 ;
        RECT 3.195 1.555 3.315 2.21 ;
        RECT 2.335 1.52 2.595 1.67 ;
        RECT 2.355 1.52 2.475 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.8 0.18 ;
        RECT 2.105 0.475 2.345 0.595 ;
        RECT 2.225 -0.18 2.345 0.595 ;
        RECT 0.685 -0.18 0.805 0.82 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.8 2.79 ;
        RECT 5.295 1.56 5.415 2.79 ;
        RECT 4.455 1.795 4.575 2.79 ;
        RECT 3.615 1.795 3.735 2.79 ;
        RECT 2.775 1.795 2.895 2.79 ;
        RECT 1.935 1.56 2.055 2.79 ;
        RECT 0.625 1.825 0.745 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.615 0.655 5.495 0.655 5.495 0.485 4.775 0.485 4.775 0.655 4.655 0.655 4.655 0.485 3.935 0.485 3.935 0.655 3.815 0.655 3.815 0.365 5.615 0.365 ;
      POLYGON 4.355 0.895 3.185 0.895 3.185 0.885 3.005 0.885 3.005 0.605 3.125 0.605 3.125 0.765 3.305 0.765 3.305 0.775 4.235 0.775 4.235 0.605 4.355 0.605 ;
      POLYGON 3.545 0.655 3.425 0.655 3.425 0.485 2.765 0.485 2.765 0.595 2.66 0.595 2.66 0.835 1.865 0.835 1.865 0.845 1.745 0.845 1.745 0.605 1.865 0.605 1.865 0.715 2.54 0.715 2.54 0.595 2.525 0.595 2.525 0.475 2.63 0.475 2.63 0.365 3.545 0.365 ;
      POLYGON 3.065 1.125 1.505 1.125 1.505 0.48 1.045 0.48 1.045 1.06 0.185 1.06 0.185 1.705 0.325 1.705 0.325 1.945 0.205 1.945 0.205 1.825 0.065 1.825 0.065 0.72 0.205 0.72 0.205 0.6 0.325 0.6 0.325 0.94 0.925 0.94 0.925 0.36 1.625 0.36 1.625 1.005 3.065 1.005 ;
      POLYGON 2.275 1.365 1.385 1.365 1.385 1.945 1.165 1.945 1.165 2.065 1.045 2.065 1.045 1.825 1.265 1.825 1.265 0.84 1.165 0.84 1.165 0.6 1.285 0.6 1.285 0.72 1.385 0.72 1.385 1.245 2.275 1.245 ;
  END
END NAND4BBX2

MACRO SDFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSXL 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.585 0.36 5.705 0.6 ;
        RECT 4.84 0.46 5.705 0.58 ;
        RECT 3.78 0.42 4.96 0.48 ;
        RECT 4.575 0.46 5.705 0.54 ;
        RECT 3.78 0.36 4.695 0.48 ;
        RECT 3.78 0.36 3.9 1.34 ;
        RECT 3.635 1.22 3.9 1.34 ;
        RECT 3.495 1.23 3.755 1.38 ;
        RECT 3.08 1.23 3.755 1.35 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.275 0.97 8.595 1.115 ;
        RECT 8.135 0.91 8.395 1.09 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.715 0.87 8.975 1.1 ;
        RECT 8.755 0.87 8.875 1.28 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.075 1.21 10.195 1.62 ;
        RECT 9.875 1.23 10.195 1.46 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.395 0.97 10.595 1.09 ;
        RECT 10.165 0.94 10.425 1.09 ;
        RECT 9.835 0.87 9.955 1.11 ;
        RECT 9.235 1.49 9.515 1.61 ;
        RECT 9.395 0.97 9.515 1.61 ;
    END
  END SE
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1644 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 0.885 1.09 1.145 ;
        RECT 0.815 0.74 0.995 1.145 ;
        RECT 0.815 0.74 0.935 2.135 ;
        RECT 0.755 0.74 0.995 0.86 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1644 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.99 0.74 2.23 0.86 ;
        RECT 1.99 0.74 2.11 1.505 ;
        RECT 1.81 1.465 2.015 1.625 ;
        RECT 1.84 1.385 2.11 1.505 ;
        RECT 1.81 1.465 1.96 1.725 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 10.315 -0.18 10.435 0.75 ;
        RECT 8.755 -0.18 8.875 0.75 ;
        RECT 6.565 -0.18 6.685 0.65 ;
        RECT 5.185 -0.18 5.425 0.34 ;
        RECT 2.92 -0.18 3.04 0.71 ;
        RECT 1.51 -0.18 1.63 0.4 ;
        RECT 0.155 0.74 0.395 0.86 ;
        RECT 0.155 -0.18 0.275 0.86 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 10.195 1.98 10.315 2.79 ;
        RECT 8.755 1.97 8.875 2.79 ;
        RECT 6.665 2.11 6.785 2.79 ;
        RECT 5.645 2.29 5.885 2.79 ;
        RECT 3.395 2.03 3.635 2.15 ;
        RECT 3.395 2.03 3.515 2.79 ;
        RECT 2.615 1.97 2.735 2.79 ;
        RECT 1.475 1.505 1.595 2.79 ;
        RECT 0.395 1.97 0.515 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.855 0.75 10.835 0.75 10.835 1.97 10.795 1.97 10.795 2.09 10.675 2.09 10.675 1.86 9.635 1.86 9.635 1.53 9.755 1.53 9.755 1.74 10.715 1.74 10.715 0.63 10.735 0.63 10.735 0.51 10.855 0.51 ;
      POLYGON 9.795 0.75 9.275 0.75 9.275 1.37 9.115 1.37 9.115 1.73 9.515 1.73 9.515 2.09 9.395 2.09 9.395 1.85 7.895 1.85 7.895 1.69 7.845 1.69 7.845 1.57 7.895 1.57 7.895 0.72 7.825 0.72 7.825 0.6 8.065 0.6 8.065 0.72 8.015 0.72 8.015 1.57 8.085 1.57 8.085 1.73 8.995 1.73 8.995 1.25 9.155 1.25 9.155 0.63 9.675 0.63 9.675 0.51 9.795 0.51 ;
      POLYGON 8.515 2.09 7.325 2.09 7.325 2.21 7.205 2.21 7.205 2.09 7.035 2.09 7.035 1.99 6.36 1.99 6.36 2.17 5.325 2.17 5.325 2.05 6.24 2.05 6.24 1.87 7.155 1.87 7.155 1.97 7.605 1.97 7.605 1.12 7.585 1.12 7.585 0.36 8.395 0.36 8.395 0.75 8.275 0.75 8.275 0.48 7.705 0.48 7.705 0.88 7.765 0.88 7.765 1.12 7.725 1.12 7.725 1.97 8.515 1.97 ;
      POLYGON 7.485 1.75 7.365 1.75 7.365 1.37 6.385 1.37 6.385 1.25 7.345 1.25 7.345 0.54 7.465 0.54 7.465 1.25 7.485 1.25 ;
      POLYGON 7.225 1.12 7.105 1.12 7.105 0.89 6.325 0.89 6.325 0.56 5.945 0.56 5.945 1.02 5.405 1.02 5.405 1.69 5.165 1.69 5.165 1.57 5.285 1.57 5.285 1.02 4.62 1.02 4.62 1.16 4.5 1.16 4.5 0.9 4.78 0.9 4.78 0.74 5.02 0.74 5.02 0.9 5.825 0.9 5.825 0.44 6.445 0.44 6.445 0.77 7.225 0.77 ;
      POLYGON 6.965 1.13 6.205 1.13 6.205 1.51 6.305 1.51 6.305 1.75 5.775 1.75 5.775 1.93 4.835 1.93 4.835 1.4 4.26 1.4 4.26 0.66 4.62 0.66 4.62 0.78 4.38 0.78 4.38 1.28 4.955 1.28 4.955 1.81 5.655 1.81 5.655 1.63 6.085 1.63 6.085 0.68 6.205 0.68 6.205 1.01 6.965 1.01 ;
      POLYGON 4.535 1.82 4.415 1.82 4.415 1.64 2.7 1.64 2.7 1.07 2.82 1.07 2.82 1.52 4.02 1.52 4.02 0.6 4.14 0.6 4.14 1.52 4.535 1.52 ;
      POLYGON 4.175 1.88 4.055 1.88 4.055 1.91 3.26 1.91 3.26 2.03 2.975 2.03 2.975 1.91 3.14 1.91 3.14 1.79 3.935 1.79 3.935 1.76 4.175 1.76 ;
      POLYGON 3.66 1.1 3.42 1.1 3.42 0.95 2.56 0.95 2.56 1.85 2.375 1.85 2.375 2.075 2.135 2.075 2.135 1.73 2.44 1.73 2.44 0.62 1.87 0.62 1.87 1.18 1.63 1.18 1.63 1.06 1.75 1.06 1.75 0.5 2.56 0.5 2.56 0.83 3.54 0.83 3.54 0.98 3.66 0.98 ;
      POLYGON 1.33 1.385 1.175 1.385 1.175 1.625 1.055 1.625 1.055 1.265 1.21 1.265 1.21 0.62 0.635 0.62 0.635 1 0.655 1 0.655 1.24 0.515 1.24 0.515 0.5 1.33 0.5 ;
  END
END SDFFSXL

MACRO MX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X4 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 1.2 1.2 1.32 ;
        RECT 0.36 1.6 1.04 1.72 ;
        RECT 0.92 1.2 1.04 1.72 ;
        RECT 0.36 1.175 0.51 1.72 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.025 0.8 1.48 ;
        RECT 0.68 1 0.8 1.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.23 2.33 1.395 ;
        RECT 1.86 1.275 2.19 1.405 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.24 1.44 3.36 2.21 ;
        RECT 3.22 0.59 3.34 0.83 ;
        RECT 3.06 1.44 3.36 1.56 ;
        RECT 3.04 0.71 3.34 0.83 ;
        RECT 2.56 1.32 3.18 1.44 ;
        RECT 2.56 0.76 3.16 0.88 ;
        RECT 2.56 1.175 2.83 1.44 ;
        RECT 2.4 1.515 2.68 1.635 ;
        RECT 2.56 0.65 2.68 1.635 ;
        RECT 2.32 0.65 2.68 0.77 ;
        RECT 2.4 1.515 2.52 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.64 -0.18 3.76 0.64 ;
        RECT 2.8 -0.18 2.92 0.64 ;
        RECT 1.9 0.46 2.14 0.58 ;
        RECT 1.9 -0.18 2.02 0.58 ;
        RECT 0.68 -0.18 0.8 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 3.66 1.56 3.78 2.79 ;
        RECT 2.82 1.56 2.94 2.79 ;
        RECT 1.98 1.56 2.1 2.79 ;
        RECT 0.64 1.84 0.76 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.44 1.11 1.74 1.11 1.74 1.84 1.4 1.84 1.4 2.21 1.28 2.21 1.28 1.72 1.62 1.72 1.62 1.11 1.56 1.11 1.56 0.64 1.32 0.64 1.32 0.4 1.44 0.4 1.44 0.52 1.68 0.52 1.68 0.99 2.44 0.99 ;
      POLYGON 1.5 1.6 1.38 1.6 1.38 1.35 1.32 1.35 1.32 1 1.12 1 1.12 0.88 0.24 0.88 0.24 1.84 0.32 1.84 0.32 2.08 0.2 2.08 0.2 1.96 0.12 1.96 0.12 0.64 0.2 0.64 0.2 0.5 0.32 0.5 0.32 0.76 1.44 0.76 1.44 1.23 1.5 1.23 ;
  END
END MX2X4

MACRO NOR4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BXL 0 0 ;
  SIZE 2.61 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.035 0.535 1.435 ;
        RECT 0.415 1.025 0.535 1.435 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 1.095 1.215 1.285 ;
        RECT 0.885 1.165 1.145 1.38 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.435 ;
        RECT 1.355 1.175 1.67 1.295 ;
        RECT 1.355 1.055 1.475 1.295 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.16 2.305 1.38 ;
        RECT 2.115 1.025 2.235 1.41 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2544 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.455 0.485 1.695 0.605 ;
        RECT 1.455 0.485 1.575 0.905 ;
        RECT 0.12 0.785 1.575 0.905 ;
        RECT 0.675 0.425 0.795 0.905 ;
        RECT 0.555 1.555 0.675 1.795 ;
        RECT 0.12 1.555 0.675 1.675 ;
        RECT 0.12 0.785 0.24 1.675 ;
        RECT 0.07 0.885 0.24 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.61 0.18 ;
        RECT 1.935 -0.18 2.055 0.665 ;
        RECT 1.095 -0.18 1.215 0.665 ;
        RECT 0.255 -0.18 0.375 0.665 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.61 2.79 ;
        RECT 1.835 1.555 1.955 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.545 1.65 2.375 1.65 2.375 1.77 2.255 1.77 2.255 1.53 2.425 1.53 2.425 0.905 1.895 0.905 1.895 1.025 1.775 1.025 1.775 0.785 2.355 0.785 2.355 0.425 2.475 0.425 2.475 0.665 2.545 0.665 ;
  END
END NOR4BXL

MACRO MXI4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X1 0 0 ;
  SIZE 6.96 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.465 0.44 2.585 1.04 ;
        RECT 2.445 0.92 2.565 1.53 ;
        RECT 1.82 0.44 2.585 0.56 ;
        RECT 1.965 0.36 2.205 0.56 ;
        RECT 0.775 0.48 1.94 0.6 ;
        RECT 0.775 0.48 0.895 1.24 ;
        RECT 0.65 0.595 0.895 0.855 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.975 1.265 3.425 1.39 ;
        RECT 2.915 1.23 3.345 1.385 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.075 1.52 4.525 1.67 ;
        RECT 4.405 1.43 4.525 1.67 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.645 1.48 4.96 1.705 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.815 1.525 6.205 1.705 ;
        RECT 5.815 1.5 6.075 1.705 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.156 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.8667 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.745 1.24 6.545 1.36 ;
        RECT 6.105 1.23 6.365 1.38 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.66 0.255 2.06 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.96 0.18 ;
        RECT 6.225 -0.18 6.345 0.38 ;
        RECT 4.825 -0.18 4.945 0.83 ;
        RECT 3.105 -0.18 3.225 0.86 ;
        RECT 1.405 -0.18 1.645 0.36 ;
        RECT 0.555 -0.18 0.795 0.32 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.96 2.79 ;
        RECT 6.145 1.94 6.265 2.79 ;
        RECT 4.54 2.065 4.66 2.79 ;
        RECT 4.42 2.065 4.66 2.185 ;
        RECT 2.985 2.22 3.225 2.79 ;
        RECT 1.225 1.91 1.465 2.03 ;
        RECT 1.225 1.91 1.345 2.79 ;
        RECT 0.495 1.88 0.735 2 ;
        RECT 0.495 1.88 0.615 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.825 0.9 6.785 0.9 6.785 1.6 6.685 1.6 6.685 2.06 6.565 2.06 6.565 1.48 6.665 1.48 6.665 0.78 6.705 0.78 6.705 0.62 5.91 0.62 5.91 0.58 5.345 0.58 5.345 0.95 5.385 0.95 5.385 1.74 5.265 1.74 5.265 1.07 4.39 1.07 4.39 0.56 3.705 0.56 3.705 1.62 3.585 1.62 3.585 0.44 4.005 0.44 4.005 0.36 4.245 0.36 4.245 0.44 4.51 0.44 4.51 0.95 5.225 0.95 5.225 0.46 5.625 0.46 5.625 0.36 5.865 0.36 5.865 0.46 6.03 0.46 6.03 0.5 6.825 0.5 ;
      POLYGON 5.705 0.82 5.625 0.82 5.625 2.06 5.505 2.06 5.505 1.98 4.975 1.98 4.975 1.945 4.3 1.945 4.3 2.25 3.385 2.25 3.385 2.1 2.865 2.1 2.865 2.25 2.625 2.25 2.625 2.13 2.745 2.13 2.745 1.98 3.505 1.98 3.505 2.13 4.18 2.13 4.18 1.825 5.095 1.825 5.095 1.86 5.505 1.86 5.505 0.82 5.465 0.82 5.465 0.7 5.705 0.7 ;
      POLYGON 5.145 1.36 4.905 1.36 4.905 1.31 4.185 1.31 4.185 1.38 4.065 1.38 4.065 1.14 4.185 1.14 4.185 1.19 5.145 1.19 ;
      POLYGON 4.105 0.8 3.945 0.8 3.945 1.89 3.865 1.89 3.865 2.01 3.745 2.01 3.745 1.86 2.625 1.86 2.625 1.99 2.505 1.99 2.505 2.11 1.825 2.11 1.825 2.25 1.585 2.25 1.585 2.13 1.705 2.13 1.705 1.99 2.385 1.99 2.385 1.87 2.505 1.87 2.505 1.74 3.825 1.74 3.825 0.68 4.105 0.68 ;
      POLYGON 2.345 0.8 2.325 0.8 2.325 1.75 2.265 1.75 2.265 1.87 2.145 1.87 2.145 1.76 0.415 1.76 0.415 1.02 0.535 1.02 0.535 1.64 2.145 1.64 2.145 1.63 2.205 1.63 2.205 0.8 2.105 0.8 2.105 0.68 2.345 0.68 ;
      POLYGON 2.085 1.51 1.215 1.51 1.215 1.52 0.975 1.52 0.975 1.4 1.095 1.4 1.095 0.84 1.015 0.84 1.015 0.72 1.255 0.72 1.255 0.84 1.215 0.84 1.215 1.39 1.965 1.39 1.965 1.27 2.085 1.27 ;
  END
END MXI4X1

MACRO OAI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.36 1.025 2.54 1.435 ;
        RECT 2.36 1.005 2.48 1.44 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.435 ;
        RECT 0.48 1.06 1.64 1.18 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.68 1.3 1.08 1.42 ;
        RECT 0.65 1.465 0.8 1.725 ;
        RECT 0.68 1.3 0.8 1.725 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.12 0.765 2.42 0.885 ;
        RECT 2.3 0.645 2.42 0.885 ;
        RECT 1.04 1.555 2.24 1.675 ;
        RECT 2.12 0.765 2.24 1.675 ;
        RECT 2.1 1.555 2.22 2.21 ;
        RECT 1.81 1.315 2.24 1.435 ;
        RECT 1.81 1.175 1.96 1.435 ;
        RECT 1.04 1.555 1.16 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 1.46 -0.18 1.58 0.7 ;
        RECT 0.62 -0.18 0.74 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.52 1.56 2.64 2.79 ;
        RECT 1.68 1.795 1.8 2.79 ;
        RECT 0.4 1.56 0.52 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.84 0.7 2.72 0.7 2.72 0.525 2 0.525 2 0.94 0.2 0.94 0.2 0.65 0.32 0.65 0.32 0.82 1.04 0.82 1.04 0.65 1.16 0.65 1.16 0.82 1.88 0.82 1.88 0.405 2.84 0.405 ;
  END
END OAI21X2

MACRO NAND4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX4 0 0 ;
  SIZE 8.41 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.035 1.08 7.635 1.2 ;
        RECT 7.035 1.08 7.275 1.35 ;
        RECT 6.675 1.26 7.235 1.38 ;
        RECT 6.975 1.23 7.275 1.35 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.315 1.08 6.555 1.2 ;
        RECT 4.945 1.26 6.435 1.38 ;
        RECT 6.315 1.08 6.435 1.38 ;
        RECT 6.105 1.23 6.435 1.38 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.265 1.26 3.845 1.38 ;
        RECT 3.495 1.23 3.755 1.38 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 1 0.395 1.24 ;
        RECT 0.07 1 0.395 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.9392 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.075 0.84 7.835 0.96 ;
        RECT 7.715 0.64 7.835 0.96 ;
        RECT 7.245 1.5 7.365 2.21 ;
        RECT 1.365 1.5 7.365 1.62 ;
        RECT 6.875 0.64 6.995 0.96 ;
        RECT 6.405 1.5 6.525 2.21 ;
        RECT 3.025 0.99 6.195 1.11 ;
        RECT 6.075 0.84 6.195 1.11 ;
        RECT 5.565 1.5 5.685 2.21 ;
        RECT 4.725 1.5 4.845 2.21 ;
        RECT 3.885 1.5 4.005 2.21 ;
        RECT 3.045 1.5 3.165 2.21 ;
        RECT 2.97 1.465 3.145 1.725 ;
        RECT 3.025 0.99 3.145 1.725 ;
        RECT 2.205 1.5 2.325 2.21 ;
        RECT 1.365 1.5 1.485 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.41 0.18 ;
        RECT 2.205 -0.18 2.325 0.69 ;
        RECT 1.365 -0.18 1.485 0.69 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.41 2.79 ;
        RECT 7.665 1.56 7.785 2.79 ;
        RECT 6.825 1.74 6.945 2.79 ;
        RECT 5.985 1.74 6.105 2.79 ;
        RECT 5.145 1.74 5.265 2.79 ;
        RECT 4.305 1.74 4.425 2.79 ;
        RECT 3.465 1.74 3.585 2.79 ;
        RECT 2.625 1.74 2.745 2.79 ;
        RECT 1.785 1.74 1.905 2.79 ;
        RECT 0.945 1.56 1.065 2.79 ;
        RECT 0.135 1.36 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.255 0.69 8.135 0.69 8.135 0.48 7.415 0.48 7.415 0.69 7.295 0.69 7.295 0.48 6.575 0.48 6.575 0.69 6.455 0.69 6.455 0.48 5.715 0.48 5.715 0.63 5.475 0.63 5.475 0.48 4.875 0.48 4.875 0.63 4.635 0.63 4.635 0.51 4.755 0.51 4.755 0.36 8.255 0.36 ;
      POLYGON 6.215 0.72 5.955 0.72 5.955 0.87 3.165 0.87 3.165 0.82 2.985 0.82 2.985 0.7 3.285 0.7 3.285 0.75 3.885 0.75 3.885 0.63 4.005 0.63 4.005 0.75 5.115 0.75 5.115 0.63 5.235 0.63 5.235 0.75 5.835 0.75 5.835 0.6 6.215 0.6 ;
      POLYGON 4.485 0.63 4.245 0.63 4.245 0.51 3.645 0.51 3.645 0.63 3.405 0.63 3.405 0.51 2.745 0.51 2.745 0.93 0.945 0.93 0.945 0.64 1.065 0.64 1.065 0.81 1.785 0.81 1.785 0.64 1.905 0.64 1.905 0.81 2.625 0.81 2.625 0.39 4.365 0.39 4.365 0.51 4.485 0.51 ;
      POLYGON 2.125 1.36 0.675 1.36 0.675 2.01 0.555 2.01 0.555 0.68 0.675 0.68 0.675 1.24 2.125 1.24 ;
  END
END NAND4BX4

MACRO TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI 0 0 ;
  SIZE 0.87 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.182 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 1.38 0.255 2.03 ;
        RECT 0.07 1.465 0.255 1.725 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 0.87 0.18 ;
        RECT 0.555 -0.18 0.675 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 0.87 2.79 ;
        RECT 0.555 1.38 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.415 1.26 0.295 1.26 0.295 0.92 0.135 0.92 0.135 0.68 0.255 0.68 0.255 0.8 0.415 0.8 ;
  END
END TIEHI

MACRO OA21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X4 0 0 ;
  SIZE 3.77 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.175 1.67 1.435 ;
        RECT 1.305 1.175 1.67 1.34 ;
        RECT 1.305 1.1 1.425 1.34 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.135 1.145 1.38 ;
        RECT 0.825 1.09 1.065 1.31 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 1.09 0.51 1.575 ;
        RECT 0.36 1.09 0.51 1.545 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.135 1.175 3.41 1.435 ;
        RECT 2.03 1.32 3.255 1.44 ;
        RECT 3.135 0.71 3.255 1.44 ;
        RECT 3.095 0.59 3.215 0.88 ;
        RECT 2.255 0.76 3.255 0.88 ;
        RECT 2.87 1.32 2.99 2.21 ;
        RECT 2.255 0.59 2.375 0.88 ;
        RECT 2.03 1.32 2.15 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.77 0.18 ;
        RECT 3.515 -0.18 3.635 0.64 ;
        RECT 2.675 -0.18 2.795 0.64 ;
        RECT 1.775 -0.18 1.895 0.53 ;
        RECT 0.625 -0.18 0.745 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.77 2.79 ;
        RECT 3.29 1.56 3.41 2.79 ;
        RECT 2.45 1.56 2.57 2.79 ;
        RECT 1.61 1.795 1.73 2.79 ;
        RECT 0.405 1.695 0.525 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.015 1.19 1.91 1.19 1.91 1.675 1.165 1.675 1.165 2.21 1.045 2.21 1.045 1.555 1.79 1.555 1.79 0.98 1.465 0.98 1.465 0.68 1.585 0.68 1.585 0.86 1.91 0.86 1.91 1.07 3.015 1.07 ;
      POLYGON 1.165 0.97 0.205 0.97 0.205 0.68 0.325 0.68 0.325 0.85 1.045 0.85 1.045 0.68 1.165 0.68 ;
  END
END OA21X4

MACRO AOI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221XL 0 0 ;
  SIZE 2.9 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 0.745 0.975 0.935 ;
        RECT 0.595 0.65 0.855 0.865 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.205 1.08 2.325 1.395 ;
        RECT 2.045 1.23 2.305 1.42 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 1.11 0.565 1.38 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 0.94 2.015 1.11 ;
        RECT 1.805 0.94 1.925 1.325 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.175 0.975 1.635 1.12 ;
        RECT 1.175 0.94 1.435 1.12 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3288 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 1.175 2.83 1.435 ;
        RECT 2.565 0.7 2.685 1.66 ;
        RECT 1.305 0.7 2.685 0.82 ;
        RECT 2.365 0.4 2.485 0.82 ;
        RECT 1.305 0.4 1.425 0.82 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.9 0.18 ;
        RECT 1.885 0.46 2.125 0.58 ;
        RECT 1.885 -0.18 2.005 0.58 ;
        RECT 0.315 -0.18 0.435 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.9 2.79 ;
        RECT 1.015 1.93 1.135 2.79 ;
        RECT 0.135 2.23 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.265 1.925 1.325 1.925 1.325 1.6 1.205 1.6 1.205 1.48 1.445 1.48 1.445 1.805 2.145 1.805 2.145 1.54 2.265 1.54 ;
      POLYGON 1.845 1.685 1.725 1.685 1.725 1.565 1.565 1.565 1.565 1.36 0.805 1.36 0.805 1.62 0.655 1.62 0.655 1.83 0.535 1.83 0.535 1.5 0.685 1.5 0.685 1.24 1.685 1.24 1.685 1.445 1.845 1.445 ;
  END
END AOI221XL

MACRO DLY2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X1 0 0 ;
  SIZE 5.51 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.82 2.54 1.145 ;
        RECT 2.33 0.94 2.45 1.26 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 1.6 0.34 2.18 ;
        RECT 0.22 0.4 0.34 0.64 ;
        RECT 0.1 0.52 0.22 1.72 ;
        RECT 0.07 1.175 0.22 1.435 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.51 0.18 ;
        RECT 4.91 1.48 5.21 1.72 ;
        RECT 5.09 0.98 5.21 1.72 ;
        RECT 4.99 -0.18 5.11 1.1 ;
        RECT 4.39 0.68 4.63 0.8 ;
        RECT 4.39 -0.18 4.51 0.8 ;
        RECT 3.19 -0.18 3.31 0.78 ;
        RECT 3.11 0.66 3.23 1.46 ;
        RECT 2.47 -0.18 2.71 0.32 ;
        RECT 1.28 1.04 1.56 1.28 ;
        RECT 1.44 -0.18 1.56 1.28 ;
        RECT 0.64 -0.18 0.76 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.51 2.79 ;
        RECT 3.91 1.22 4.97 1.34 ;
        RECT 4.29 1.92 4.53 2.79 ;
        RECT 4.29 1.7 4.41 2.79 ;
        RECT 3.91 1.7 4.41 1.82 ;
        RECT 3.91 1 4.03 1.82 ;
        RECT 2.49 2.18 2.73 2.3 ;
        RECT 2.495 2.18 2.615 2.79 ;
        RECT 1.08 0.76 1.32 0.9 ;
        RECT 0.34 0.76 1.32 0.88 ;
        RECT 0.46 1.88 0.76 2.79 ;
        RECT 0.46 1.36 0.58 2.79 ;
        RECT 0.34 0.76 0.46 1.48 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 5.45 1.98 4.99 1.98 4.99 1.96 4.67 1.96 4.67 1.58 4.15 1.58 4.15 1.46 4.79 1.46 4.79 1.84 5.33 1.84 5.33 0.86 5.23 0.86 5.23 0.62 5.35 0.62 5.35 0.74 5.45 0.74 ;
      POLYGON 4.87 1.04 4.15 1.04 4.15 0.5 3.55 0.5 3.55 1.7 3.37 1.7 3.37 1.82 3.25 1.82 3.25 1.58 3.43 1.58 3.43 0.38 4.27 0.38 4.27 0.92 4.75 0.92 4.75 0.48 4.63 0.48 4.63 0.36 4.87 0.36 ;
      POLYGON 4.17 2.06 2.37 2.06 2.37 2.25 0.925 2.25 0.925 1.88 0.88 1.88 0.88 1.76 0.7 1.76 0.7 1.24 0.58 1.24 0.58 1 0.7 1 0.7 1.12 0.82 1.12 0.82 1.64 1 1.64 1 1.76 1.045 1.76 1.045 2.13 2.25 2.13 2.25 1.94 3.67 1.94 3.67 0.76 3.91 0.76 3.91 0.62 4.03 0.62 4.03 0.88 3.79 0.88 3.79 1.94 4.17 1.94 ;
      POLYGON 3.07 0.54 2.95 0.54 2.95 0.56 1.8 0.56 1.8 1.52 1.54 1.52 1.54 1.77 1.42 1.77 1.42 1.4 1.68 1.4 1.68 0.4 1.8 0.4 1.8 0.44 2.83 0.44 2.83 0.42 3.07 0.42 ;
      POLYGON 2.19 1.82 2.13 1.82 2.13 2.01 1.18 2.01 1.18 1.64 1.12 1.64 1.12 1.52 0.94 1.52 0.94 1.19 1.06 1.19 1.06 1.4 1.24 1.4 1.24 1.52 1.3 1.52 1.3 1.89 2.01 1.89 2.01 1.7 2.07 1.7 2.07 0.68 2.19 0.68 ;
  END
END DLY2X1

MACRO OAI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X4 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.79 0.97 4.295 1.09 ;
        RECT 3.79 0.82 3.91 1.09 ;
        RECT 2.2 0.82 3.91 0.94 ;
        RECT 1.855 0.97 2.32 1.09 ;
        RECT 2.045 0.94 2.32 1.09 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.095 1.09 5.215 1.33 ;
        RECT 5 0.885 5.15 1.21 ;
        RECT 4.565 1.09 5.215 1.21 ;
        RECT 3.34 1.21 4.685 1.33 ;
        RECT 3.34 1.06 3.46 1.33 ;
        RECT 2.545 1.06 3.46 1.18 ;
        RECT 1.525 1.21 2.665 1.33 ;
        RECT 2.545 1.06 2.665 1.33 ;
        RECT 1.525 0.99 1.645 1.33 ;
        RECT 0.875 0.99 1.645 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.93 1.45 5.555 1.57 ;
        RECT 5.435 1.24 5.555 1.57 ;
        RECT 2.785 1.3 3.025 1.57 ;
        RECT 0.93 1.32 1.05 1.57 ;
        RECT 0.595 1.32 1.05 1.44 ;
        RECT 0.595 1.23 0.855 1.44 ;
        RECT 0.595 1.2 0.715 1.44 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.375 1.225 7.075 1.345 ;
        RECT 6.685 1.225 6.945 1.38 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.1072 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.095 0.65 7.335 0.77 ;
        RECT 6.135 0.76 7.215 0.88 ;
        RECT 6.915 1.56 7.035 2.21 ;
        RECT 1.835 1.69 7.035 1.81 ;
        RECT 6.135 0.65 6.495 0.88 ;
        RECT 6.135 1.465 6.31 1.81 ;
        RECT 6.135 0.65 6.255 1.81 ;
        RECT 6.075 1.56 6.195 2.21 ;
        RECT 4.395 1.69 4.515 2.21 ;
        RECT 1.835 1.69 1.955 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 5.355 0.34 5.595 0.46 ;
        RECT 5.355 -0.18 5.475 0.46 ;
        RECT 4.395 0.34 4.635 0.46 ;
        RECT 4.395 -0.18 4.515 0.46 ;
        RECT 3.435 0.34 3.675 0.46 ;
        RECT 3.435 -0.18 3.555 0.46 ;
        RECT 2.475 0.34 2.715 0.46 ;
        RECT 2.475 -0.18 2.595 0.46 ;
        RECT 1.515 0.34 1.755 0.46 ;
        RECT 1.515 -0.18 1.635 0.46 ;
        RECT 0.555 0.34 0.795 0.46 ;
        RECT 0.555 -0.18 0.675 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.335 1.56 7.455 2.79 ;
        RECT 6.495 1.93 6.615 2.79 ;
        RECT 5.655 1.93 5.775 2.79 ;
        RECT 3.015 1.93 3.135 2.79 ;
        RECT 0.455 1.56 0.575 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.695 0.65 7.575 0.65 7.575 0.53 6.855 0.53 6.855 0.64 6.735 0.64 6.735 0.53 6.015 0.53 6.015 0.7 0.075 0.7 0.075 0.58 5.895 0.58 5.895 0.41 6.735 0.41 6.735 0.4 6.855 0.4 6.855 0.41 7.695 0.41 ;
  END
END OAI31X4

MACRO TLATNTSCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX12 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.305 0.82 0.565 1.09 ;
        RECT 0.305 0.78 0.545 1.09 ;
    END
  END E
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 0.76 1.09 1.205 ;
        RECT 0.925 0.78 1.045 1.25 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 0.76 1.385 1.25 ;
        RECT 1.23 0.76 1.385 1.22 ;
    END
  END CK
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.925 1.31 11.045 2.21 ;
        RECT 10.085 1.04 11.045 1.16 ;
        RECT 10.925 0.405 11.045 1.16 ;
        RECT 10.745 1.31 11.045 1.43 ;
        RECT 7.585 1.19 10.865 1.31 ;
        RECT 10.085 1.04 10.865 1.31 ;
        RECT 10.085 0.405 10.205 2.21 ;
        RECT 9.245 0.405 9.365 2.21 ;
        RECT 8.405 1.04 9.365 1.31 ;
        RECT 8.405 0.405 8.525 2.21 ;
        RECT 7.585 1.175 7.76 1.435 ;
        RECT 7.585 0.8 7.705 1.45 ;
        RECT 7.565 1.33 7.685 2.21 ;
        RECT 7.565 0.4 7.685 0.92 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 11.345 -0.18 11.465 0.92 ;
        RECT 10.505 -0.18 10.625 0.92 ;
        RECT 9.665 -0.18 9.785 0.92 ;
        RECT 8.825 -0.18 8.945 0.92 ;
        RECT 7.985 -0.18 8.105 0.92 ;
        RECT 7.145 -0.18 7.265 0.64 ;
        RECT 6.045 0.47 6.285 0.59 ;
        RECT 6.045 -0.18 6.165 0.59 ;
        RECT 4.765 -0.18 4.885 0.58 ;
        RECT 2.935 0.69 3.175 0.81 ;
        RECT 2.935 -0.18 3.055 0.81 ;
        RECT 1.065 -0.18 1.185 0.64 ;
        RECT 0.225 -0.18 0.345 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 11.345 1.43 11.465 2.79 ;
        RECT 10.505 1.43 10.625 2.79 ;
        RECT 9.665 1.43 9.785 2.79 ;
        RECT 8.825 1.43 8.945 2.79 ;
        RECT 7.985 1.43 8.105 2.79 ;
        RECT 7.085 1.72 7.325 2.15 ;
        RECT 7.085 1.72 7.205 2.79 ;
        RECT 6.305 1.72 6.425 2.79 ;
        RECT 5.465 1.72 5.585 2.79 ;
        RECT 4.625 1.44 4.745 2.79 ;
        RECT 3.295 2.13 3.415 2.79 ;
        RECT 3.175 2.13 3.415 2.25 ;
        RECT 1.005 1.61 1.125 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.465 1.21 7.085 1.21 7.085 1.6 6.845 1.6 6.845 2.21 6.725 2.21 6.725 1.6 6.005 1.6 6.005 2.21 5.885 2.21 5.885 1.6 5.165 1.6 5.165 2.09 5.045 2.09 5.045 1.48 6.965 1.48 6.965 0.88 6.745 0.88 6.745 0.83 5.525 0.83 5.525 0.78 5.405 0.78 5.405 0.66 5.645 0.66 5.645 0.71 6.745 0.71 6.745 0.6 6.865 0.6 6.865 0.76 7.085 0.76 7.085 1.09 7.465 1.09 ;
      POLYGON 6.845 1.12 5.165 1.12 5.165 0.82 4.525 0.82 4.525 0.48 3.775 0.48 3.775 0.76 3.735 0.76 3.735 1.29 3.075 1.29 3.075 1.65 3.895 1.65 3.895 1.89 4.015 1.89 4.015 2.01 3.775 2.01 3.775 1.77 2.955 1.77 2.955 1.37 2.835 1.37 2.835 1.17 3.615 1.17 3.615 0.64 3.655 0.64 3.655 0.36 4.645 0.36 4.645 0.7 5.285 0.7 5.285 1 6.845 1 ;
      POLYGON 6.225 1.36 4.925 1.36 4.925 1.06 4.265 1.06 4.265 1.68 4.145 1.68 4.145 1.53 3.195 1.53 3.195 1.41 4.145 1.41 4.145 0.72 4.285 0.72 4.285 0.6 4.405 0.6 4.405 0.94 5.045 0.94 5.045 1.24 6.225 1.24 ;
      POLYGON 4.625 1.3 4.505 1.3 4.505 1.92 4.45 1.92 4.45 2.25 3.535 2.25 3.535 2.01 2.655 2.01 2.655 2.11 2.535 2.11 2.535 1.99 2.355 1.99 2.355 0.82 2.235 0.82 2.235 0.7 2.475 0.7 2.475 1.87 2.655 1.87 2.655 1.89 3.655 1.89 3.655 2.13 4.33 2.13 4.33 1.8 4.385 1.8 4.385 1.18 4.625 1.18 ;
      POLYGON 3.535 0.48 3.415 0.48 3.415 1.05 2.715 1.05 2.715 1.51 2.795 1.51 2.795 1.75 2.675 1.75 2.675 1.63 2.595 1.63 2.595 0.58 2.33 0.58 2.33 0.52 1.625 0.52 1.625 1.49 1.605 1.49 1.605 1.73 1.485 1.73 1.485 1.37 1.505 1.37 1.505 0.64 1.485 0.64 1.485 0.4 2.095 0.4 2.095 0.38 2.335 0.38 2.335 0.4 2.45 0.4 2.45 0.46 2.815 0.46 2.815 0.93 3.295 0.93 3.295 0.36 3.535 0.36 ;
      POLYGON 2.235 2.07 2.115 2.07 2.115 1.97 1.245 1.97 1.245 1.49 0.485 1.49 0.485 1.73 0.365 1.73 0.365 1.37 0.685 1.37 0.685 0.66 0.645 0.66 0.645 0.4 0.765 0.4 0.765 0.54 0.805 0.54 0.805 1.37 1.365 1.37 1.365 1.85 1.935 1.85 1.935 0.82 1.815 0.82 1.815 0.7 2.055 0.7 2.055 1.83 2.235 1.83 ;
  END
END TLATNTSCAX12

MACRO NAND3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BXL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.04 0.51 1.51 ;
        RECT 0.36 1.04 0.48 1.54 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.81 1.02 0.935 1.26 ;
        RECT 0.65 1.02 0.935 1.145 ;
        RECT 0.65 0.885 0.805 1.145 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.515 1.355 1.67 1.735 ;
        RECT 1.48 1.355 1.67 1.725 ;
    END
  END AN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.915 1.84 1.155 1.96 ;
        RECT 0.915 1.66 1.035 1.96 ;
        RECT 0.12 1.66 1.035 1.78 ;
        RECT 0.12 0.8 0.455 0.92 ;
        RECT 0.335 0.68 0.455 0.92 ;
        RECT 0.135 1.66 0.255 2.02 ;
        RECT 0.07 1.465 0.24 1.725 ;
        RECT 0.12 0.8 0.24 1.78 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.295 -0.18 1.415 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.395 1.9 1.515 2.79 ;
        RECT 0.555 1.9 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.935 2.02 1.815 2.02 1.815 1.9 1.79 1.9 1.79 1.235 1.15 1.235 1.15 1.115 1.715 1.115 1.715 0.68 1.835 0.68 1.835 0.995 1.91 0.995 1.91 1.78 1.935 1.78 ;
  END
END NAND3BXL

MACRO CLKINVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX12 0 0 ;
  SIZE 4.64 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.296 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.755 1.15 3.835 1.27 ;
        RECT 0.885 1.15 1.145 1.38 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.0736 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 1.5 4.075 1.62 ;
        RECT 3.955 0.91 4.075 1.62 ;
        RECT 3.915 1.43 4.035 2.21 ;
        RECT 0.555 0.91 4.075 1.03 ;
        RECT 3.915 0.4 4.035 1.03 ;
        RECT 3.84 1.465 4.035 1.725 ;
        RECT 3.075 1.43 3.195 2.21 ;
        RECT 3.075 0.4 3.195 1.03 ;
        RECT 2.235 1.43 2.355 2.21 ;
        RECT 2.235 0.4 2.355 1.03 ;
        RECT 1.395 1.43 1.515 2.21 ;
        RECT 1.395 0.4 1.515 1.03 ;
        RECT 0.555 1.43 0.675 2.21 ;
        RECT 0.555 0.4 0.675 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.64 0.18 ;
        RECT 4.335 -0.18 4.455 0.915 ;
        RECT 3.495 -0.18 3.615 0.79 ;
        RECT 2.655 -0.18 2.775 0.79 ;
        RECT 1.815 -0.18 1.935 0.79 ;
        RECT 0.975 -0.18 1.095 0.79 ;
        RECT 0.135 -0.18 0.255 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.64 2.79 ;
        RECT 4.335 1.43 4.455 2.79 ;
        RECT 3.495 1.74 3.615 2.79 ;
        RECT 2.655 1.74 2.775 2.79 ;
        RECT 1.815 1.74 1.935 2.79 ;
        RECT 0.975 1.74 1.095 2.79 ;
        RECT 0.135 1.43 0.255 2.79 ;
    END
  END VDD
END CLKINVX12

MACRO OAI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X1 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.09 0.785 2.25 1.215 ;
        RECT 2.09 0.77 2.21 1.215 ;
    END
  END B0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.03 2.85 1.435 ;
        RECT 2.73 1.015 2.85 1.435 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.115 1.09 1.435 ;
        RECT 0.86 1.01 0.98 1.32 ;
    END
  END A1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 0.77 2.54 1.22 ;
        RECT 2.41 0.77 2.53 1.26 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.04 0.51 1.495 ;
        RECT 0.39 1.01 0.51 1.495 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.52 1.03 1.69 1.435 ;
        RECT 1.57 1.015 1.69 1.435 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7811 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 1.465 3.12 1.725 ;
        RECT 2.97 0.775 3.09 1.725 ;
        RECT 2.89 1.555 3.01 2.21 ;
        RECT 2.67 0.775 3.09 0.895 ;
        RECT 1.41 1.555 3.12 1.675 ;
        RECT 2.67 0.6 2.79 0.895 ;
        RECT 1.41 1.555 1.53 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 1.02 -0.18 1.14 0.65 ;
        RECT 0.18 -0.18 0.3 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.25 1.795 2.37 2.79 ;
        RECT 0.38 1.615 0.5 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.21 0.65 3.09 0.65 3.09 0.53 2.91 0.53 2.91 0.48 2.37 0.48 2.37 0.65 2.25 0.65 2.25 0.48 1.53 0.48 1.53 0.65 1.41 0.65 1.41 0.36 3.03 0.36 3.03 0.41 3.21 0.41 ;
      POLYGON 1.95 0.89 0.6 0.89 0.6 0.6 0.72 0.6 0.72 0.77 1.83 0.77 1.83 0.6 1.95 0.6 ;
  END
END OAI222X1

MACRO CLKMX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X4 0 0 ;
  SIZE 4.06 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.146 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.92 1.2 1.2 1.32 ;
        RECT 0.36 1.6 1.04 1.72 ;
        RECT 0.92 1.2 1.04 1.72 ;
        RECT 0.36 1.175 0.51 1.72 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.025 0.8 1.48 ;
        RECT 0.68 1 0.8 1.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.045 1.23 2.33 1.395 ;
        RECT 1.86 1.275 2.19 1.405 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.24 1.44 3.36 2.21 ;
        RECT 3.22 0.59 3.34 0.83 ;
        RECT 3.06 1.44 3.36 1.56 ;
        RECT 3.04 0.71 3.34 0.83 ;
        RECT 2.56 1.32 3.18 1.44 ;
        RECT 2.56 0.76 3.16 0.88 ;
        RECT 2.56 1.175 2.83 1.44 ;
        RECT 2.4 1.515 2.68 1.635 ;
        RECT 2.56 0.65 2.68 1.635 ;
        RECT 2.32 0.65 2.68 0.77 ;
        RECT 2.4 1.515 2.52 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.06 0.18 ;
        RECT 3.64 -0.18 3.76 0.64 ;
        RECT 2.8 -0.18 2.92 0.64 ;
        RECT 1.9 0.46 2.14 0.58 ;
        RECT 1.9 -0.18 2.02 0.58 ;
        RECT 0.68 -0.18 0.8 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.06 2.79 ;
        RECT 3.66 1.56 3.78 2.79 ;
        RECT 2.82 1.56 2.94 2.79 ;
        RECT 1.98 1.56 2.1 2.79 ;
        RECT 0.64 1.84 0.76 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.44 1.11 1.74 1.11 1.74 1.84 1.4 1.84 1.4 2.21 1.28 2.21 1.28 1.72 1.62 1.72 1.62 1.11 1.56 1.11 1.56 0.64 1.32 0.64 1.32 0.4 1.44 0.4 1.44 0.52 1.68 0.52 1.68 0.99 2.44 0.99 ;
      POLYGON 1.5 1.6 1.38 1.6 1.38 1.35 1.32 1.35 1.32 1 1.12 1 1.12 0.88 0.24 0.88 0.24 1.84 0.32 1.84 0.32 2.08 0.2 2.08 0.2 1.96 0.12 1.96 0.12 0.64 0.2 0.64 0.2 0.5 0.32 0.5 0.32 0.76 1.44 0.76 1.44 1.23 1.5 1.23 ;
  END
END CLKMX2X4

MACRO EDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX2 0 0 ;
  SIZE 13.34 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.175 0.645 1.41 ;
        RECT 0.525 1.17 0.645 1.41 ;
        RECT 0.36 1.175 0.51 1.435 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.015 1.25 2.405 1.37 ;
        RECT 1.025 1.81 2.135 1.93 ;
        RECT 2.015 1.25 2.135 1.93 ;
        RECT 1.025 1.17 1.145 1.93 ;
        RECT 0.885 1.52 1.145 1.67 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.465 1.25 4.585 1.56 ;
        RECT 4.42 1.44 4.57 1.755 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.455 1.23 10.715 1.445 ;
        RECT 10.565 0.97 10.685 1.445 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.255 1.175 11.53 1.435 ;
        RECT 11.115 1.55 11.375 1.67 ;
        RECT 11.255 0.59 11.375 1.67 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.075 1.55 12.315 1.67 ;
        RECT 12.075 1.175 12.215 1.67 ;
        RECT 12.095 0.59 12.215 1.67 ;
        RECT 11.96 1.175 12.215 1.435 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 13.34 0.18 ;
        RECT 12.515 -0.18 12.635 0.64 ;
        RECT 11.675 -0.18 11.795 0.64 ;
        RECT 10.835 -0.18 10.955 0.79 ;
        RECT 9.485 -0.18 9.725 0.38 ;
        RECT 7.585 0.53 7.825 0.65 ;
        RECT 7.585 -0.18 7.705 0.65 ;
        RECT 5.565 0.53 5.805 0.65 ;
        RECT 5.685 -0.18 5.805 0.65 ;
        RECT 4.155 -0.18 4.275 0.65 ;
        RECT 2.755 0.53 2.995 0.65 ;
        RECT 2.755 -0.18 2.875 0.65 ;
        RECT 2.425 -0.18 2.545 0.65 ;
        RECT 0.845 -0.18 0.965 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 13.34 2.79 ;
        RECT 12.615 2.15 12.735 2.79 ;
        RECT 11.595 2.03 11.835 2.15 ;
        RECT 11.595 2.03 11.715 2.79 ;
        RECT 10.695 2.09 10.815 2.79 ;
        RECT 9.425 1.68 9.665 1.81 ;
        RECT 9.425 1.68 9.545 2.79 ;
        RECT 7.585 2.29 7.825 2.79 ;
        RECT 5.625 2.15 5.745 2.79 ;
        RECT 4.445 2.21 4.565 2.79 ;
        RECT 0.785 2.29 1.025 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 13.205 1.73 13.085 1.73 13.085 1.35 12.335 1.35 12.335 1.23 12.995 1.23 12.995 0.59 13.115 0.59 13.115 1.23 13.205 1.23 ;
      POLYGON 13.055 2.19 12.935 2.19 12.935 2.03 12.73 2.03 12.73 1.91 10.82 1.91 10.82 1.97 10.025 1.97 10.025 2.16 9.905 2.16 9.905 1.56 9.305 1.56 9.305 2.21 9.185 2.21 9.185 2.17 6.21 2.17 6.21 2.03 5.27 2.03 5.27 2.05 5.005 2.05 5.005 2.09 3.945 2.09 3.945 2.25 3.825 2.25 3.825 1.97 4.885 1.97 4.885 1.93 5.15 1.93 5.15 1.91 6.33 1.91 6.33 2.05 9.165 2.05 9.165 1.44 9.905 1.44 9.905 0.74 10.205 0.74 10.205 0.86 10.025 0.86 10.025 1.85 10.7 1.85 10.7 1.79 10.875 1.79 10.875 1.29 10.975 1.29 10.975 0.91 11.095 0.91 11.095 1.41 10.995 1.41 10.995 1.79 12.85 1.79 12.85 1.91 13.055 1.91 ;
      POLYGON 10.535 0.79 10.445 0.79 10.445 1.11 10.335 1.11 10.335 1.73 10.215 1.73 10.215 0.99 10.325 0.99 10.325 0.62 9.19 0.62 9.19 0.5 8.545 0.5 8.545 1.25 8.565 1.25 8.565 1.37 8.325 1.37 8.325 1.25 8.425 1.25 8.425 0.5 8.065 0.5 8.065 0.89 7.205 0.89 7.205 1.43 7.085 1.43 7.085 0.56 6.405 0.56 6.405 1.13 5.415 1.13 5.415 1.01 6.285 1.01 6.285 0.44 7.205 0.44 7.205 0.77 7.945 0.77 7.945 0.38 8.925 0.38 8.925 0.36 9.165 0.36 9.165 0.38 9.31 0.38 9.31 0.5 10.535 0.5 ;
      POLYGON 9.745 1.24 9.625 1.24 9.625 1.08 8.805 1.08 8.805 1.69 8.565 1.69 8.565 1.57 8.685 1.57 8.685 0.84 8.845 0.84 8.845 0.62 8.965 0.62 8.965 0.96 9.745 0.96 ;
      POLYGON 9.165 1.32 9.045 1.32 9.045 1.93 6.54 1.93 6.54 1.49 6.485 1.49 6.485 1.37 5.315 1.37 5.315 1.75 5.195 1.75 5.195 1.49 5.175 1.49 5.175 1.13 4.965 1.13 4.965 0.68 5.205 0.68 5.205 1.01 5.295 1.01 5.295 1.25 6.725 1.25 6.725 1.37 6.66 1.37 6.66 1.81 8.925 1.81 8.925 1.2 9.165 1.2 ;
      POLYGON 8.305 1.13 8.205 1.13 8.205 1.57 8.305 1.57 8.305 1.69 8.065 1.69 8.065 1.57 8.085 1.57 8.085 1.13 7.605 1.13 7.605 1.14 7.365 1.14 7.365 1.02 7.485 1.02 7.485 1.01 8.185 1.01 8.185 0.62 8.305 0.62 ;
      POLYGON 7.965 1.37 7.845 1.37 7.845 1.67 7.02 1.67 7.02 1.69 6.78 1.69 6.78 1.57 6.845 1.57 6.845 0.8 6.525 0.8 6.525 0.68 6.965 0.68 6.965 1.55 7.725 1.55 7.725 1.25 7.965 1.25 ;
      POLYGON 6.165 0.48 6.045 0.48 6.045 0.89 5.325 0.89 5.325 0.56 5.19 0.56 5.19 0.5 4.515 0.5 4.515 0.89 3.795 0.89 3.795 1.13 2.855 1.13 2.855 1.75 2.735 1.75 2.735 1.13 1.895 1.13 1.895 1.69 1.655 1.69 1.655 1.57 1.775 1.57 1.775 1.01 1.725 1.01 1.725 0.6 1.845 0.6 1.845 0.89 1.895 0.89 1.895 1.01 3.675 1.01 3.675 0.62 3.795 0.62 3.795 0.74 3.985 0.74 3.985 0.77 4.395 0.77 4.395 0.38 5.31 0.38 5.31 0.44 5.445 0.44 5.445 0.77 5.925 0.77 5.925 0.36 6.165 0.36 ;
      POLYGON 4.925 1.81 4.805 1.81 4.805 1.69 4.705 1.69 4.705 1.13 4.245 1.13 4.245 1.25 4.125 1.25 4.125 1.01 4.635 1.01 4.635 0.62 4.755 0.62 4.755 0.89 4.825 0.89 4.825 1.57 4.925 1.57 ;
      POLYGON 4.085 1.81 3.965 1.81 3.965 1.57 3.245 1.57 3.245 1.81 3.125 1.81 3.125 1.45 4.085 1.45 ;
      POLYGON 3.665 2.05 2.375 2.05 2.375 1.81 2.255 1.81 2.255 1.69 2.495 1.69 2.495 1.93 3.545 1.93 3.545 1.69 3.665 1.69 ;
      POLYGON 3.355 0.48 3.235 0.48 3.235 0.89 2.055 0.89 2.055 0.48 1.385 0.48 1.385 1.57 1.505 1.57 1.505 1.69 1.265 1.69 1.265 0.36 2.175 0.36 2.175 0.77 3.115 0.77 3.115 0.36 3.355 0.36 ;
      POLYGON 2.065 2.17 0.365 2.17 0.365 1.675 0.12 1.675 0.12 0.93 0.425 0.93 0.425 0.68 0.545 0.68 0.545 1.05 0.24 1.05 0.24 1.555 0.485 1.555 0.485 2.05 2.065 2.05 ;
  END
END EDFFTRX2

MACRO OA21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X2 0 0 ;
  SIZE 3.19 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.23 0.77 1.38 1.145 ;
        RECT 1.25 0.77 1.37 1.26 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.175 0.95 1.295 ;
        RECT 0.83 1.055 0.95 1.295 ;
        RECT 0.65 1.175 0.8 1.435 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.125 0.51 1.56 ;
        RECT 0.39 1.08 0.51 1.56 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.13 0.65 2.43 0.77 ;
        RECT 1.89 1.005 2.25 1.145 ;
        RECT 2.13 0.65 2.25 1.145 ;
        RECT 2.1 0.885 2.25 1.145 ;
        RECT 1.89 1.005 2.01 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.19 0.18 ;
        RECT 2.67 -0.18 2.79 0.64 ;
        RECT 1.77 -0.18 1.89 0.53 ;
        RECT 0.615 -0.18 0.735 0.4 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.19 2.79 ;
        RECT 2.31 1.56 2.43 2.79 ;
        RECT 1.47 1.62 1.59 2.79 ;
        RECT 0.35 1.68 0.47 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.77 1.48 1.62 1.48 1.62 1.5 1.19 1.5 1.19 1.535 1.11 1.535 1.11 1.8 0.99 1.8 0.99 1.415 1.07 1.415 1.07 1.38 1.5 1.38 1.5 0.68 1.62 0.68 1.62 1.24 1.77 1.24 ;
      POLYGON 1.11 0.92 0.99 0.92 0.99 0.86 0.075 0.86 0.075 0.74 0.99 0.74 0.99 0.68 1.11 0.68 ;
  END
END OA21X2

MACRO OAI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X2 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 0.975 3.7 1.44 ;
        RECT 3.55 0.945 3.67 1.44 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.61 0.885 2.83 1.145 ;
        RECT 0.65 0.82 2.8 0.94 ;
        RECT 2.61 0.82 2.73 1.15 ;
        RECT 0.65 0.82 0.77 1.15 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.93 1.06 2.45 1.18 ;
        RECT 1.23 1.06 1.38 1.435 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.87 1.3 2.11 1.42 ;
        RECT 1.755 1.52 2.015 1.67 ;
        RECT 1.87 1.3 2.015 1.67 ;
    END
  END A2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.31 0.65 3.67 0.77 ;
        RECT 1.79 1.79 3.43 1.91 ;
        RECT 3.31 0.65 3.43 1.91 ;
        RECT 2.97 1.56 3.43 1.91 ;
        RECT 3.17 1.56 3.29 2.21 ;
        RECT 2.97 1.465 3.12 1.91 ;
        RECT 1.79 1.79 1.91 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 2.53 0.34 2.77 0.46 ;
        RECT 2.53 -0.18 2.65 0.46 ;
        RECT 1.57 0.34 1.81 0.46 ;
        RECT 1.57 -0.18 1.69 0.46 ;
        RECT 0.61 0.34 0.85 0.46 ;
        RECT 0.61 -0.18 0.73 0.46 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.59 1.56 3.71 2.79 ;
        RECT 2.69 2.03 2.93 2.15 ;
        RECT 2.69 2.03 2.81 2.79 ;
        RECT 0.51 1.56 0.63 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.03 0.65 3.91 0.65 3.91 0.53 3.19 0.53 3.19 0.7 0.13 0.7 0.13 0.58 3.07 0.58 3.07 0.41 4.03 0.41 ;
  END
END OAI31X2

MACRO EDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX4 0 0 ;
  SIZE 11.6 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.16 0.51 1.63 ;
        RECT 0.375 1.16 0.495 1.66 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.365 1.295 5.605 1.49 ;
        RECT 5.235 1.23 5.495 1.45 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.305 1.25 6.895 1.37 ;
        RECT 6.395 1.23 6.655 1.38 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.695 1.315 8.815 2.21 ;
        RECT 7.9 1.315 8.815 1.435 ;
        RECT 7.445 0.72 8.645 0.84 ;
        RECT 7.9 1.175 8.05 1.435 ;
        RECT 7.9 0.72 8.02 1.555 ;
        RECT 7.855 1.435 7.975 2.21 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.365 0.72 10.565 0.84 ;
        RECT 10.375 1.32 10.495 2.21 ;
        RECT 9.64 1.32 10.495 1.44 ;
        RECT 9.64 1.175 9.79 1.44 ;
        RECT 9.64 0.72 9.76 1.56 ;
        RECT 9.535 1.44 9.655 2.21 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.6 0.18 ;
        RECT 10.925 -0.18 11.045 0.71 ;
        RECT 9.845 -0.18 10.085 0.36 ;
        RECT 8.885 -0.18 9.125 0.36 ;
        RECT 7.925 -0.18 8.165 0.36 ;
        RECT 6.965 -0.18 7.205 0.32 ;
        RECT 5.105 -0.18 5.225 0.79 ;
        RECT 4.205 0.61 4.445 0.73 ;
        RECT 4.205 -0.18 4.325 0.73 ;
        RECT 2.545 0.61 2.785 0.73 ;
        RECT 2.545 -0.18 2.665 0.73 ;
        RECT 0.555 -0.18 0.675 0.8 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.6 2.79 ;
        RECT 10.795 1.58 10.915 2.79 ;
        RECT 9.955 1.56 10.075 2.79 ;
        RECT 9.115 1.56 9.235 2.79 ;
        RECT 8.275 1.56 8.395 2.79 ;
        RECT 7.435 1.74 7.555 2.79 ;
        RECT 5.325 2.17 5.565 2.29 ;
        RECT 5.325 2.17 5.445 2.79 ;
        RECT 4.365 2.17 4.605 2.29 ;
        RECT 4.365 2.17 4.485 2.79 ;
        RECT 2.545 1.81 2.785 1.93 ;
        RECT 2.545 1.81 2.665 2.79 ;
        RECT 0.555 1.78 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 11.465 0.9 11.335 0.9 11.335 2.21 11.215 2.21 11.215 1.46 10.615 1.46 10.615 1.22 10.735 1.22 10.735 1.34 11.215 1.34 11.215 0.78 11.345 0.78 11.345 0.66 11.465 0.66 ;
      POLYGON 11.095 1.22 10.975 1.22 10.975 0.95 10.685 0.95 10.685 0.6 8.925 0.6 8.925 1.16 8.685 1.16 8.685 1.04 8.805 1.04 8.805 0.6 6.285 0.6 6.285 0.79 6.165 0.79 6.165 0.49 5.49 0.49 5.49 1.03 4.985 1.03 4.985 1.69 5.085 1.69 5.085 1.81 4.845 1.81 4.845 1.69 4.865 1.69 4.865 1.17 4.125 1.17 4.125 1.05 4.685 1.05 4.685 0.65 4.805 0.65 4.805 0.77 4.985 0.77 4.985 0.91 5.37 0.91 5.37 0.37 6.285 0.37 6.285 0.48 10.805 0.48 10.805 0.83 11.095 0.83 ;
      POLYGON 7.695 1.62 6.685 1.62 6.685 1.87 6.565 1.87 6.565 1.5 7.575 1.5 7.575 1.24 7.695 1.24 ;
      POLYGON 7.135 1.86 7.015 1.86 7.015 1.98 6.925 1.98 6.925 2.11 6.445 2.11 6.445 2.25 5.885 2.25 5.885 2.13 6.325 2.13 6.325 1.62 6.065 1.62 6.065 1.05 5.965 1.05 5.965 0.93 6.405 0.93 6.405 0.72 6.735 0.72 6.735 0.84 6.525 0.84 6.525 1.05 6.185 1.05 6.185 1.5 6.445 1.5 6.445 1.99 6.805 1.99 6.805 1.86 6.895 1.86 6.895 1.74 7.135 1.74 ;
      POLYGON 6.205 2.01 5.41 2.01 5.41 2.05 4.085 2.05 4.085 2.11 2.905 2.11 2.905 1.69 2.425 1.69 2.425 2.11 1.51 2.11 1.51 1.99 1.485 1.99 1.485 1.75 1.305 1.75 1.305 0.76 1.365 0.76 1.365 0.64 1.485 0.64 1.485 0.88 1.425 0.88 1.425 1.63 1.605 1.63 1.605 1.87 1.63 1.87 1.63 1.99 2.305 1.99 2.305 1.57 3.025 1.57 3.025 1.99 3.965 1.99 3.965 1.93 5.29 1.93 5.29 1.89 5.725 1.89 5.725 0.73 5.685 0.73 5.685 0.61 5.925 0.61 5.925 0.73 5.845 0.73 5.845 1.74 6.205 1.74 ;
      POLYGON 4.745 1.55 4.725 1.55 4.725 1.79 3.745 1.79 3.745 1.81 3.505 1.81 3.505 1.69 3.565 1.69 3.565 0.64 3.685 0.64 3.685 1.67 4.605 1.67 4.605 1.43 4.625 1.43 4.625 1.31 4.745 1.31 ;
      POLYGON 3.985 1.55 3.865 1.55 3.865 0.52 3.025 0.52 3.025 0.97 2.305 0.97 2.305 0.52 1.725 0.52 1.725 1.37 1.785 1.37 1.785 1.49 1.545 1.49 1.545 1.37 1.605 1.37 1.605 0.52 1.195 0.52 1.195 0.56 1.095 0.56 1.095 1.9 0.975 1.9 0.975 0.44 1.075 0.44 1.075 0.4 2.005 0.4 2.005 0.36 2.245 0.36 2.245 0.4 2.425 0.4 2.425 0.85 2.905 0.85 2.905 0.4 3.345 0.4 3.345 0.36 3.585 0.36 3.585 0.4 3.985 0.4 ;
      POLYGON 3.265 1.87 3.145 1.87 3.145 1.21 2.325 1.21 2.325 1.09 3.145 1.09 3.145 0.64 3.265 0.64 ;
      POLYGON 3.005 1.45 2.085 1.45 2.085 1.75 2.025 1.75 2.025 1.87 1.905 1.87 1.905 1.63 1.965 1.63 1.965 0.82 1.845 0.82 1.845 0.7 2.085 0.7 2.085 1.33 3.005 1.33 ;
      POLYGON 0.835 1.16 0.715 1.16 0.715 1.04 0.24 1.04 0.24 1.75 0.255 1.75 0.255 1.99 0.135 1.99 0.135 1.87 0.12 1.87 0.12 0.8 0.135 0.8 0.135 0.56 0.255 0.56 0.255 0.92 0.835 0.92 ;
  END
END EDFFX4

MACRO EDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX1 0 0 ;
  SIZE 8.12 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.09 0.51 1.545 ;
        RECT 0.36 1.07 0.48 1.545 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.265 1.23 7.525 1.46 ;
        RECT 7.275 1.08 7.395 1.49 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.555 0.94 7.815 1.09 ;
        RECT 7.555 0.94 7.795 1.11 ;
        RECT 6.945 0.84 7.675 0.96 ;
        RECT 7.105 0.36 7.225 0.96 ;
        RECT 6.345 0.36 7.225 0.48 ;
        RECT 6.945 0.84 7.065 1.15 ;
        RECT 6.345 0.36 6.465 1.46 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.085 1.53 5.405 1.65 ;
        RECT 5.085 0.63 5.205 1.65 ;
        RECT 5 1.175 5.205 1.435 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 8.12 0.18 ;
        RECT 7.445 -0.18 7.565 0.72 ;
        RECT 5.565 -0.18 5.685 0.73 ;
        RECT 4.485 0.5 4.725 0.62 ;
        RECT 4.485 -0.18 4.605 0.62 ;
        RECT 2.705 0.43 2.945 0.55 ;
        RECT 2.705 -0.18 2.825 0.55 ;
        RECT 0.555 -0.18 0.675 0.71 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 8.12 2.79 ;
        RECT 7.385 1.85 7.505 2.79 ;
        RECT 5.625 2.1 5.865 2.22 ;
        RECT 5.625 2.1 5.745 2.79 ;
        RECT 4.685 2.01 4.925 2.13 ;
        RECT 4.685 2.01 4.805 2.79 ;
        RECT 2.795 1.75 2.915 2.79 ;
        RECT 0.555 1.665 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 8.055 1.73 7.985 1.73 7.985 1.85 7.865 1.85 7.865 1.73 6.945 1.73 6.945 1.42 6.825 1.42 6.825 1.3 7.065 1.3 7.065 1.61 7.935 1.61 7.935 0.72 7.865 0.72 7.865 0.48 7.985 0.48 7.985 0.6 8.055 0.6 ;
      POLYGON 6.985 0.72 6.705 0.72 6.705 1.56 6.765 1.56 6.765 2.21 6.645 2.21 6.645 1.98 5.85 1.98 5.85 1.89 4.38 1.89 4.38 2.23 3.085 2.23 3.085 1.63 2.675 1.63 2.675 2.23 1.525 2.23 1.525 1.59 1.365 1.59 1.365 0.72 1.305 0.72 1.305 0.6 1.545 0.6 1.545 0.72 1.485 0.72 1.485 1.47 1.645 1.47 1.645 2.11 2.555 2.11 2.555 1.51 3.205 1.51 3.205 2.11 4.26 2.11 4.26 1.77 5.97 1.77 5.97 1.86 6.645 1.86 6.645 1.68 6.585 1.68 6.585 0.6 6.985 0.6 ;
      POLYGON 6.405 1.74 6.09 1.74 6.09 1.41 5.505 1.41 5.505 1.29 6.09 1.29 6.09 0.77 5.985 0.77 5.985 0.65 6.225 0.65 6.225 0.77 6.21 0.77 6.21 1.62 6.405 1.62 ;
      POLYGON 5.965 1.09 5.725 1.09 5.725 0.97 5.325 0.97 5.325 0.51 4.965 0.51 4.965 0.86 4.545 0.86 4.545 1.63 4.065 1.63 4.065 1.99 3.945 1.99 3.945 1.47 4.065 1.47 4.065 1.51 4.425 1.51 4.425 0.86 3.925 0.86 3.925 0.78 3.905 0.78 3.905 0.54 4.025 0.54 4.025 0.66 4.045 0.66 4.045 0.74 4.845 0.74 4.845 0.39 5.445 0.39 5.445 0.85 5.845 0.85 5.845 0.97 5.965 0.97 ;
      POLYGON 4.305 1.39 4.185 1.39 4.185 1.1 3.665 1.1 3.665 1.06 3.565 1.06 3.565 0.94 3.665 0.94 3.665 0.48 3.185 0.48 3.185 0.79 2.385 0.79 2.385 1.12 2.225 1.12 2.225 0.88 2.265 0.88 2.265 0.48 1.785 0.48 1.785 1.21 1.845 1.21 1.845 1.33 1.605 1.33 1.605 1.21 1.665 1.21 1.665 0.48 1.135 0.48 1.135 1.665 1.095 1.665 1.095 1.785 0.975 1.785 0.975 1.545 1.015 1.545 1.015 0.71 0.975 0.71 0.975 0.36 2.585 0.36 2.585 0.67 3.065 0.67 3.065 0.36 3.785 0.36 3.785 0.94 3.805 0.94 3.805 0.98 4.305 0.98 ;
      POLYGON 3.545 0.72 3.445 0.72 3.445 1.99 3.325 1.99 3.325 1.39 2.745 1.39 2.745 1.15 2.865 1.15 2.865 1.27 3.325 1.27 3.325 0.72 3.305 0.72 3.305 0.6 3.545 0.6 ;
      POLYGON 3.205 1.15 3.085 1.15 3.085 1.03 2.625 1.03 2.625 1.36 2.105 1.36 2.105 1.99 1.985 1.99 1.985 0.72 1.905 0.72 1.905 0.6 2.145 0.6 2.145 0.72 2.105 0.72 2.105 1.24 2.505 1.24 2.505 0.91 3.205 0.91 ;
      POLYGON 0.895 0.99 0.655 0.99 0.655 0.95 0.24 0.95 0.24 1.665 0.255 1.665 0.255 1.905 0.135 1.905 0.135 1.785 0.12 1.785 0.12 0.71 0.135 0.71 0.135 0.47 0.255 0.47 0.255 0.83 0.895 0.83 ;
  END
END EDFFHQX1

MACRO SDFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX2 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.245 1.09 1.38 1.525 ;
        RECT 1.215 1.09 1.38 1.505 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.172 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.565 1.22 2.885 1.41 ;
        RECT 2.565 1.18 2.805 1.41 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.645 0.93 7.765 1.17 ;
        RECT 7.32 0.93 7.765 1.05 ;
        RECT 7.32 0.885 7.47 1.145 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.965 1.255 9.265 1.485 ;
        RECT 9.005 1.23 9.265 1.485 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.005 0.99 9.525 1.11 ;
        RECT 8.125 0.97 9.265 1.09 ;
        RECT 8.715 0.94 8.975 1.09 ;
        RECT 8.125 0.97 8.245 1.44 ;
    END
  END SE
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.585 1.465 0.8 1.725 ;
        RECT 0.575 1.38 0.77 1.5 ;
        RECT 0.585 1.38 0.705 2.03 ;
        RECT 0.575 0.8 0.695 1.5 ;
        RECT 0.555 0.68 0.675 0.92 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.185 -0.18 9.305 0.82 ;
        RECT 7.645 -0.18 7.765 0.64 ;
        RECT 4.985 -0.18 5.225 0.39 ;
        RECT 2.705 0.38 2.945 0.5 ;
        RECT 2.705 -0.18 2.825 0.5 ;
        RECT 0.975 -0.18 1.095 0.73 ;
        RECT 0.135 -0.18 0.255 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 9.025 1.845 9.145 2.79 ;
        RECT 7.525 2.28 7.765 2.79 ;
        RECT 5.585 2.26 5.825 2.79 ;
        RECT 4.745 2.01 4.865 2.79 ;
        RECT 4.625 2.01 4.865 2.13 ;
        RECT 3.005 2.01 3.125 2.79 ;
        RECT 2.885 2.01 3.125 2.13 ;
        RECT 1.985 2.01 2.105 2.79 ;
        RECT 1.005 1.625 1.125 2.79 ;
        RECT 0.165 1.38 0.285 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.765 1.725 9.625 1.725 9.625 1.845 9.505 1.845 9.505 1.725 8.525 1.725 8.525 1.24 8.645 1.24 8.645 1.605 9.645 1.605 9.645 0.82 9.605 0.82 9.605 0.58 9.725 0.58 9.725 0.7 9.765 0.7 ;
      POLYGON 8.665 0.82 8.005 0.82 8.005 1.56 8.405 1.56 8.405 2.21 8.285 2.21 8.285 1.68 8.005 1.68 8.005 1.8 7.74 1.8 7.74 1.98 6.835 1.98 6.835 1.3 6.445 1.3 6.445 0.6 6.745 0.6 6.745 0.72 6.565 0.72 6.565 1.18 6.955 1.18 6.955 1.86 7.62 1.86 7.62 1.68 7.885 1.68 7.885 0.7 8.545 0.7 8.545 0.56 8.665 0.56 ;
      POLYGON 7.405 1.74 7.08 1.74 7.08 1.06 6.685 1.06 6.685 0.94 6.865 0.94 6.865 0.48 5.965 0.48 5.965 0.86 6.085 0.86 6.085 1.1 5.845 1.1 5.845 0.63 4.745 0.63 4.745 0.48 4.265 0.48 4.265 0.99 4.445 0.99 4.445 1.11 4.145 1.11 4.145 0.36 4.865 0.36 4.865 0.51 5.845 0.51 5.845 0.36 6.985 0.36 6.985 0.59 7.2 0.59 7.2 1.62 7.405 1.62 ;
      POLYGON 7.405 2.22 5.945 2.22 5.945 2.14 5.25 2.14 5.25 2.01 4.985 2.01 4.985 1.89 4.29 1.89 4.29 2.23 3.325 2.23 3.325 1.89 1.425 1.89 1.425 1.645 1.5 1.645 1.5 0.92 1.455 0.92 1.455 0.68 1.575 0.68 1.575 0.8 1.62 0.8 1.62 1.77 3.325 1.77 3.325 0.86 3.445 0.86 3.445 2.11 3.905 2.11 3.905 1.15 4.025 1.15 4.025 2.11 4.17 2.11 4.17 1.77 5.105 1.77 5.105 1.89 5.37 1.89 5.37 2.02 6.065 2.02 6.065 2.1 7.405 2.1 ;
      POLYGON 6.535 1.94 6.415 1.94 6.415 1.54 6.205 1.54 6.205 1.34 4.925 1.34 4.925 1.11 4.805 1.11 4.805 0.99 5.045 0.99 5.045 1.22 6.205 1.22 6.205 0.72 6.085 0.72 6.085 0.6 6.325 0.6 6.325 1.42 6.535 1.42 ;
      POLYGON 6.115 1.9 5.995 1.9 5.995 1.78 5.73 1.78 5.73 1.77 5.225 1.77 5.225 1.65 5.105 1.65 5.105 1.53 5.345 1.53 5.345 1.65 5.85 1.65 5.85 1.66 6.115 1.66 ;
      POLYGON 5.725 1.1 5.605 1.1 5.605 0.87 4.685 0.87 4.685 1.65 4.145 1.65 4.145 1.53 4.565 1.53 4.565 0.87 4.385 0.87 4.385 0.6 4.625 0.6 4.625 0.75 5.725 0.75 ;
      POLYGON 3.785 1.99 3.665 1.99 3.665 0.74 2.205 0.74 2.205 1.12 2.085 1.12 2.085 0.62 3.665 0.62 3.665 0.54 3.785 0.54 ;
      POLYGON 3.085 1.1 2.965 1.1 2.965 1.06 2.445 1.06 2.445 1.53 2.645 1.53 2.645 1.65 2.325 1.65 2.325 1.36 1.845 1.36 1.845 0.56 1.335 0.56 1.335 0.97 0.935 0.97 0.935 1.26 0.815 1.26 0.815 0.85 1.215 0.85 1.215 0.44 1.965 0.44 1.965 1.24 2.325 1.24 2.325 0.94 2.965 0.94 2.965 0.86 3.085 0.86 ;
  END
END SDFFRHQX2

MACRO SDFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX2 0 0 ;
  SIZE 15.08 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.575 0.36 1.695 1.7 ;
        RECT 0.895 0.36 1.695 0.48 ;
        RECT 0.975 0.94 1.215 1.06 ;
        RECT 0.39 0.9 1.095 1.02 ;
        RECT 0.895 0.36 1.015 1.02 ;
        RECT 0.36 1.175 0.51 1.435 ;
        RECT 0.39 0.9 0.51 1.435 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.735 1.14 0.855 1.57 ;
        RECT 0.65 1.14 0.855 1.555 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.885 2.25 1.145 ;
        RECT 1.815 0.9 2.25 1.02 ;
        RECT 1.815 0.9 1.935 1.14 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.39 1.035 2.54 1.5 ;
        RECT 2.39 0.96 2.51 1.5 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.876 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.3 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.945 0.945 5.33 1.12 ;
        RECT 4.945 0.94 5.205 1.14 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.195 1.12 12.455 1.38 ;
        RECT 12.185 1.1 12.425 1.34 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.905 0.68 13.025 2.03 ;
        RECT 12.83 1.465 13.025 1.725 ;
        RECT 12.86 1.38 13.025 1.725 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 13.725 0.74 14.045 0.86 ;
        RECT 13.745 1.3 13.865 2.03 ;
        RECT 13.725 0.74 13.845 1.42 ;
        RECT 13.41 1.025 13.845 1.145 ;
        RECT 13.41 0.885 13.56 1.145 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 15.08 0.18 ;
        RECT 14.285 -0.18 14.525 0.32 ;
        RECT 13.325 -0.18 13.565 0.32 ;
        RECT 12.365 -0.18 12.605 0.32 ;
        RECT 11.21 -0.18 11.33 0.83 ;
        RECT 4.99 -0.18 5.23 0.32 ;
        RECT 2.9 -0.18 3.02 0.92 ;
        RECT 1.86 -0.18 1.98 0.78 ;
        RECT 0.555 -0.18 0.675 0.78 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 15.08 2.79 ;
        RECT 14.165 1.38 14.285 2.79 ;
        RECT 13.325 1.38 13.445 2.79 ;
        RECT 12.485 1.5 12.605 2.79 ;
        RECT 10.95 2.13 11.07 2.79 ;
        RECT 10.83 2.13 11.07 2.25 ;
        RECT 8.45 1.88 8.57 2.79 ;
        RECT 8.33 1.88 8.57 2 ;
        RECT 6.23 1.96 6.35 2.79 ;
        RECT 6.11 1.96 6.35 2.08 ;
        RECT 4.85 2.13 4.97 2.79 ;
        RECT 2.925 2.28 3.165 2.79 ;
        RECT 2.055 1.86 2.175 2.79 ;
        RECT 0.695 1.93 0.815 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 15.005 0.86 14.885 0.86 14.885 1.18 14.705 1.18 14.705 1.62 14.585 1.62 14.585 1.18 13.965 1.18 13.965 1.06 14.765 1.06 14.765 0.74 15.005 0.74 ;
      POLYGON 14.885 0.52 14.765 0.52 14.765 0.56 13.265 0.56 13.265 1.26 13.145 1.26 13.145 0.56 12.785 0.56 12.785 1.26 12.665 1.26 12.665 0.6 11.75 0.6 11.75 0.84 11.71 0.84 11.71 1.59 11.55 1.59 11.55 2.01 11.43 2.01 11.43 1.47 11.59 1.47 11.59 1.11 10.49 1.11 10.49 0.99 11.59 0.99 11.59 0.72 11.63 0.72 11.63 0.48 12.665 0.48 12.665 0.44 14.645 0.44 14.645 0.4 14.885 0.4 ;
      POLYGON 12.2 0.84 12.065 0.84 12.065 1.62 12.185 1.62 12.185 2.25 11.19 2.25 11.19 2.01 8.93 2.01 8.93 1.52 8.11 1.52 8.11 1.4 9.05 1.4 9.05 1.89 11.31 1.89 11.31 2.13 12.065 2.13 12.065 1.74 11.945 1.74 11.945 0.72 12.2 0.72 ;
      POLYGON 11.47 1.35 9.41 1.35 9.41 1.04 7.61 1.04 7.61 1.6 7.55 1.6 7.55 1.72 7.43 1.72 7.43 1.48 7.49 1.48 7.49 0.62 7.61 0.62 7.61 0.92 9.53 0.92 9.53 1.23 11.47 1.23 ;
      POLYGON 10.91 0.83 10.79 0.83 10.79 0.59 10.67 0.59 10.67 0.53 10.13 0.53 10.13 0.77 9.89 0.77 9.89 0.65 10.01 0.65 10.01 0.41 10.79 0.41 10.79 0.47 10.91 0.47 ;
      POLYGON 10.71 2.25 8.69 2.25 8.69 1.76 8.21 1.76 8.21 1.96 7.68 1.96 7.68 2.2 6.47 2.2 6.47 1.84 5.99 1.84 5.99 2.25 5.11 2.25 5.11 2.13 5.87 2.13 5.87 1.72 6.59 1.72 6.59 2.08 7.56 2.08 7.56 1.84 8.09 1.84 8.09 1.64 8.81 1.64 8.81 2.13 10.71 2.13 ;
      POLYGON 10.59 1.77 9.17 1.77 9.17 1.28 7.99 1.28 7.99 1.52 7.97 1.52 7.97 1.72 7.85 1.72 7.85 1.4 7.87 1.4 7.87 1.16 9.29 1.16 9.29 1.65 10.59 1.65 ;
      POLYGON 10.55 0.77 10.37 0.77 10.37 1.01 9.65 1.01 9.65 0.8 7.85 0.8 7.85 0.68 9.77 0.68 9.77 0.89 10.25 0.89 10.25 0.65 10.55 0.65 ;
      POLYGON 7.81 0.48 7.37 0.48 7.37 1.28 7.31 1.28 7.31 1.96 6.71 1.96 6.71 1.6 5.75 1.6 5.75 2.01 4.96 2.01 4.96 1.62 4.43 1.62 4.43 1.14 4.55 1.14 4.55 1.5 5.08 1.5 5.08 1.89 5.63 1.89 5.63 1.48 6.83 1.48 6.83 1.84 7.19 1.84 7.19 1.16 7.25 1.16 7.25 0.36 7.81 0.36 ;
      POLYGON 7.13 1.04 7.07 1.04 7.07 1.72 6.95 1.72 6.95 1.36 5.445 1.36 5.445 1.65 5.51 1.65 5.51 1.77 5.27 1.77 5.27 1.65 5.325 1.65 5.325 1.38 4.73 1.38 4.73 1.26 5.325 1.26 5.325 1.24 6.17 1.24 6.17 0.62 6.29 0.62 6.29 1.24 6.95 1.24 6.95 0.92 7.01 0.92 7.01 0.62 7.13 0.62 ;
      POLYGON 6.71 0.86 6.59 0.86 6.59 0.74 6.46 0.74 6.46 0.5 6.05 0.5 6.05 0.8 5.69 0.8 5.69 0.68 5.93 0.68 5.93 0.38 6.58 0.38 6.58 0.62 6.71 0.62 ;
      POLYGON 5.81 0.48 5.69 0.48 5.69 0.56 4.75 0.56 4.75 0.5 4.07 0.5 4.07 1.63 4.03 1.63 4.03 1.75 3.91 1.75 3.91 1.51 3.95 1.51 3.95 0.5 3.44 0.5 3.44 0.8 3.55 0.8 3.55 1.7 3.54 1.7 3.54 1.82 3.42 1.82 3.42 1.58 3.43 1.58 3.43 0.92 3.32 0.92 3.32 0.38 4.365 0.38 4.365 0.36 4.605 0.36 4.605 0.38 4.87 0.38 4.87 0.44 5.57 0.44 5.57 0.36 5.81 0.36 ;
      POLYGON 5.79 1.12 5.45 1.12 5.45 0.82 4.31 0.82 4.31 1.97 4.27 1.97 4.27 2.09 4.15 2.09 4.15 1.85 4.19 1.85 4.19 0.68 4.43 0.68 4.43 0.7 5.57 0.7 5.57 1 5.79 1 ;
      POLYGON 3.85 2.21 3.73 2.21 3.73 2.16 2.295 2.16 2.295 1.74 1.935 1.74 1.935 1.94 1.455 1.94 1.455 2.05 1.335 2.05 1.335 0.72 1.135 0.72 1.135 0.6 1.455 0.6 1.455 1.82 1.815 1.82 1.815 1.62 2.415 1.62 2.415 2.04 3.67 2.04 3.67 0.74 3.71 0.74 3.71 0.62 3.83 0.62 3.83 0.86 3.79 0.86 3.79 1.97 3.85 1.97 ;
      POLYGON 3.31 1.42 2.78 1.42 2.78 1.92 2.535 1.92 2.535 1.8 2.66 1.8 2.66 0.72 2.255 0.72 2.255 0.6 2.78 0.6 2.78 1.3 3.31 1.3 ;
      POLYGON 1.195 1.81 0.375 1.81 0.375 2.05 0.255 2.05 0.255 1.93 0.12 1.93 0.12 0.935 0.135 0.935 0.135 0.54 0.255 0.54 0.255 1.055 0.24 1.055 0.24 1.69 1.075 1.69 1.075 1.22 1.195 1.22 ;
  END
END SDFFSRX2

MACRO NAND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4XL 0 0 ;
  SIZE 2.03 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 1.025 1.535 1.265 ;
        RECT 1.23 1.025 1.535 1.145 ;
        RECT 1.23 0.885 1.38 1.145 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 0.88 1.11 1.285 ;
        RECT 0.94 0.75 1.09 1.145 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.595 0.8 1.045 ;
        RECT 0.67 0.595 0.79 1.245 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.595 0.51 1.015 ;
        RECT 0.35 0.805 0.47 1.245 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2976 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 1.405 1.775 1.525 ;
        RECT 1.655 0.785 1.775 1.525 ;
        RECT 1.52 0.665 1.675 0.855 ;
        RECT 1.52 0.595 1.67 0.855 ;
        RECT 1.55 0.785 1.775 0.905 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.03 0.18 ;
        RECT 0.135 -0.18 0.255 0.385 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.03 2.79 ;
        RECT 1.775 1.985 1.895 2.79 ;
        RECT 0.855 1.985 0.975 2.79 ;
        RECT 0.135 1.985 0.255 2.79 ;
    END
  END VDD
END NAND4XL

MACRO CLKAND2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X3 0 0 ;
  SIZE 3.48 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.151 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.265 1.02 1.665 1.14 ;
        RECT 0.595 0.97 1.385 1.09 ;
        RECT 0.595 0.94 0.855 1.09 ;
        RECT 0.435 1.02 0.765 1.14 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.151 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 1.21 1.145 1.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.648 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.225 1.25 3.345 2.14 ;
        RECT 2.39 1.25 3.345 1.37 ;
        RECT 2.265 0.79 3.045 0.91 ;
        RECT 2.925 0.62 3.045 0.91 ;
        RECT 2.39 0.79 2.54 1.37 ;
        RECT 2.385 1.27 2.51 1.39 ;
        RECT 2.385 1.27 2.505 2.14 ;
        RECT 2.025 0.68 2.385 0.8 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 3.48 0.18 ;
        RECT 2.505 -0.18 2.625 0.67 ;
        RECT 1.605 0.49 1.845 0.61 ;
        RECT 1.605 -0.18 1.725 0.61 ;
        RECT 0.335 -0.18 0.455 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 3.48 2.79 ;
        RECT 2.805 1.49 2.925 2.79 ;
        RECT 1.905 2.095 2.025 2.79 ;
        RECT 1.035 2.095 1.155 2.79 ;
        RECT 0.135 1.575 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.27 1.15 1.905 1.15 1.905 1.72 0.495 1.72 0.495 1.6 1.785 1.6 1.785 0.85 1.065 0.85 1.065 0.8 0.945 0.8 0.945 0.68 1.185 0.68 1.185 0.73 1.905 0.73 1.905 1.03 2.27 1.03 ;
  END
END CLKAND2X3

MACRO EDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX2 0 0 ;
  SIZE 9.86 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 1.15 0.855 1.38 ;
        RECT 0.605 1.12 0.725 1.53 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.375 1.075 6.615 1.28 ;
        RECT 6.45 1.075 6.6 1.47 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.975 1.23 7.235 1.38 ;
        RECT 5.835 1.83 7.15 1.95 ;
        RECT 7.03 1.14 7.15 1.95 ;
        RECT 6.99 1.14 7.15 1.38 ;
        RECT 5.515 1.99 5.955 2.11 ;
        RECT 5.835 1.39 5.955 2.11 ;
        RECT 5.775 0.92 5.895 1.51 ;
        RECT 5.655 0.92 5.895 1.04 ;
        RECT 5.395 2.13 5.635 2.25 ;
        RECT 5.515 1.99 5.635 2.25 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.73 0.94 8.105 1.09 ;
        RECT 7.73 0.74 7.865 1.09 ;
        RECT 7.73 0.74 7.85 1.65 ;
        RECT 7.69 1.53 7.81 2.18 ;
        RECT 7.625 0.74 7.865 0.86 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.51 0.74 8.825 0.86 ;
        RECT 8.53 1.53 8.65 2.18 ;
        RECT 8.51 0.74 8.63 1.65 ;
        RECT 8.48 0.885 8.63 1.145 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.86 0.18 ;
        RECT 9.065 -0.18 9.305 0.38 ;
        RECT 8.165 -0.18 8.285 0.38 ;
        RECT 7.145 -0.18 7.385 0.38 ;
        RECT 6.235 -0.18 6.475 0.38 ;
        RECT 4.695 -0.18 4.815 0.73 ;
        RECT 2.815 -0.18 3.055 0.32 ;
        RECT 0.705 0.58 0.945 0.7 ;
        RECT 0.705 -0.18 0.825 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.86 2.79 ;
        RECT 8.95 1.53 9.07 2.79 ;
        RECT 8.11 1.57 8.23 2.79 ;
        RECT 7.27 1.53 7.39 2.79 ;
        RECT 6.235 2.07 6.475 2.19 ;
        RECT 6.235 2.07 6.355 2.79 ;
        RECT 4.575 1.97 4.815 2.09 ;
        RECT 4.575 1.97 4.695 2.79 ;
        RECT 2.815 2.26 3.055 2.79 ;
        RECT 0.765 1.65 0.885 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.785 0.86 9.665 0.86 9.665 1.31 9.55 1.31 9.55 1.77 9.43 1.77 9.43 1.31 8.75 1.31 8.75 1.19 9.545 1.19 9.545 0.74 9.785 0.74 ;
      POLYGON 9.665 0.54 9.545 0.54 9.545 0.62 8.345 0.62 8.345 1.45 7.97 1.45 7.97 1.21 8.225 1.21 8.225 0.62 7.505 0.62 7.505 1 7.525 1 7.525 1.24 7.385 1.24 7.385 0.62 5.895 0.62 5.895 0.48 5.235 0.48 5.235 0.97 5.215 0.97 5.215 1.49 5.295 1.49 5.295 1.61 5.055 1.61 5.055 1.49 5.095 1.49 5.095 0.97 4.695 0.97 4.695 1.12 4.375 1.12 4.375 1 4.575 1 4.575 0.85 5.115 0.85 5.115 0.36 6.015 0.36 6.015 0.5 9.425 0.5 9.425 0.42 9.665 0.42 ;
      POLYGON 6.91 1.71 6.67 1.71 6.67 1.59 6.735 1.59 6.735 0.955 6.255 0.955 6.255 1.26 6.015 1.26 6.015 0.835 6.665 0.835 6.665 0.74 6.905 0.74 6.905 0.86 6.855 0.86 6.855 1.59 6.91 1.59 ;
      POLYGON 5.775 0.72 5.535 0.72 5.535 1.63 5.715 1.63 5.715 1.87 5.595 1.87 5.595 1.85 4.39 1.85 4.39 1.9 1.735 1.9 1.735 1.66 1.575 1.66 1.575 0.8 1.515 0.8 1.515 0.68 1.755 0.68 1.755 0.8 1.695 0.8 1.695 1.54 1.855 1.54 1.855 1.78 4.27 1.78 4.27 1.73 5.415 1.73 5.415 0.6 5.775 0.6 ;
      POLYGON 4.975 1.33 4.935 1.33 4.935 1.58 4.115 1.58 4.115 1.66 3.775 1.66 3.775 0.62 3.895 0.62 3.895 1.46 4.815 1.46 4.815 1.21 4.855 1.21 4.855 1.09 4.975 1.09 ;
      POLYGON 4.255 1.34 4.015 1.34 4.015 0.5 3.55 0.5 3.55 0.56 1.995 0.56 1.995 1.22 2.055 1.22 2.055 1.34 1.815 1.34 1.815 1.22 1.875 1.22 1.875 0.56 1.325 0.56 1.325 1.65 1.305 1.65 1.305 1.77 1.185 1.77 1.185 1.53 1.205 1.53 1.205 0.76 1.185 0.76 1.185 0.44 2.255 0.44 2.255 0.36 2.495 0.36 2.495 0.44 3.43 0.44 3.43 0.38 3.575 0.38 3.575 0.36 3.815 0.36 3.815 0.38 4.135 0.38 4.135 1.22 4.255 1.22 ;
      RECT 2.275 2.02 3.855 2.14 ;
      POLYGON 3.575 1.66 3.335 1.66 3.335 1.02 2.775 1.02 2.775 1.2 2.655 1.2 2.655 0.9 3.295 0.9 3.295 0.68 3.535 0.68 3.535 0.8 3.455 0.8 3.455 1.54 3.575 1.54 ;
      POLYGON 3.215 1.44 2.335 1.44 2.335 1.66 2.095 1.66 2.095 1.54 2.215 1.54 2.215 0.8 2.115 0.8 2.115 0.68 2.355 0.68 2.355 0.8 2.335 0.8 2.335 1.32 3.095 1.32 3.095 1.14 3.215 1.14 ;
      POLYGON 1.085 1.02 0.845 1.02 0.845 1 0.465 1 0.465 1.77 0.345 1.77 0.345 0.52 0.465 0.52 0.465 0.88 1.085 0.88 ;
  END
END EDFFX2

MACRO CLKAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X6 0 0 ;
  SIZE 5.8 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.105 0.94 3.225 1.24 ;
        RECT 0.595 0.94 3.225 1.06 ;
        RECT 1.535 0.94 1.775 1.11 ;
        RECT 0.385 0.99 0.855 1.11 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.895 1.18 2.505 1.3 ;
        RECT 1.755 1.23 2.015 1.38 ;
        RECT 1.295 1.23 2.015 1.35 ;
        RECT 1.145 1.18 1.415 1.3 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.2237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.545 1.39 5.665 2.21 ;
        RECT 3.865 1.39 5.665 1.51 ;
        RECT 5.405 0.4 5.525 0.915 ;
        RECT 5.225 0.795 5.525 0.915 ;
        RECT 3.665 0.91 5.345 1.03 ;
        RECT 4.745 1.175 5.15 1.51 ;
        RECT 4.745 0.795 4.865 1.51 ;
        RECT 4.705 1.39 4.825 2.21 ;
        RECT 4.565 0.795 4.865 1.03 ;
        RECT 4.565 0.4 4.685 1.03 ;
        RECT 3.865 1.39 3.985 2.21 ;
        RECT 3.665 0.4 3.785 1.03 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 5.8 0.18 ;
        RECT 4.985 -0.18 5.105 0.79 ;
        RECT 4.145 -0.18 4.265 0.79 ;
        RECT 3.185 0.46 3.425 0.58 ;
        RECT 3.185 -0.18 3.305 0.58 ;
        RECT 1.695 0.46 1.935 0.58 ;
        RECT 1.695 -0.18 1.815 0.58 ;
        RECT 0.285 -0.18 0.405 0.64 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 5.8 2.79 ;
        RECT 5.125 1.63 5.245 2.79 ;
        RECT 4.285 1.63 4.405 2.79 ;
        RECT 3.385 2.045 3.505 2.79 ;
        RECT 2.545 2.045 2.665 2.79 ;
        RECT 1.825 2.045 1.945 2.79 ;
        RECT 0.985 2.045 1.105 2.79 ;
        RECT 0.135 2.045 0.255 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.625 1.27 3.465 1.27 3.465 1.62 0.445 1.62 0.445 1.5 3.345 1.5 3.345 0.82 1.175 0.82 1.175 0.77 1.055 0.77 1.055 0.65 1.295 0.65 1.295 0.7 2.545 0.7 2.545 0.65 2.785 0.65 2.785 0.7 3.465 0.7 3.465 1.15 4.625 1.15 ;
  END
END CLKAND2X6

MACRO DLY3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X1 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 1.465 2.925 1.725 ;
        RECT 2.705 1.405 2.925 1.725 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3024 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.365 1.23 4.625 1.38 ;
        RECT 4.405 1.11 4.525 2.21 ;
        RECT 4.265 1.11 4.525 1.23 ;
        RECT 4.265 0.68 4.385 1.23 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.11 1.48 7.53 1.72 ;
        RECT 7.41 0.98 7.53 1.72 ;
        RECT 7.205 0.98 7.53 1.1 ;
        RECT 7.205 -0.18 7.325 1.1 ;
        RECT 6.725 0.62 6.845 0.86 ;
        RECT 6.605 -0.18 6.725 0.74 ;
        RECT 5.325 1.22 5.565 1.34 ;
        RECT 5.445 -0.18 5.565 1.34 ;
        RECT 4.745 0.6 4.985 0.72 ;
        RECT 4.845 -0.18 4.965 0.72 ;
        RECT 3.635 1.465 3.875 1.585 ;
        RECT 3.635 -0.18 3.755 1.585 ;
        RECT 2.835 -0.18 2.955 0.885 ;
        RECT 1.875 0.76 1.995 1.52 ;
        RECT 1.575 0.76 1.995 0.88 ;
        RECT 1.575 -0.18 1.695 0.88 ;
        RECT 1.175 -0.18 1.295 0.64 ;
        RECT 0.375 1.32 0.795 1.44 ;
        RECT 0.375 -0.18 0.495 1.44 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 6.165 1.22 7.29 1.34 ;
        RECT 6.61 1.92 6.73 2.79 ;
        RECT 6.23 1.22 6.35 2.79 ;
        RECT 4.765 1.7 5.005 2.15 ;
        RECT 4.865 1.7 4.985 2.79 ;
        RECT 3.275 1.245 3.515 1.365 ;
        RECT 3.275 1.245 3.395 2.79 ;
        RECT 2.925 1.845 3.045 2.79 ;
        RECT 0.615 1 1.755 1.12 ;
        RECT 1.175 1.89 1.675 2.01 ;
        RECT 1.555 1 1.675 2.01 ;
        RECT 1.175 1.89 1.435 2.79 ;
        RECT 1.055 1.8 1.295 1.92 ;
        RECT 0.615 0.78 0.855 1.12 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.77 1.98 7.19 1.98 7.19 1.96 6.87 1.96 6.87 1.66 6.47 1.66 6.47 1.54 6.99 1.54 6.99 1.84 7.65 1.84 7.65 0.86 7.445 0.86 7.445 0.62 7.565 0.62 7.565 0.74 7.77 0.74 ;
      POLYGON 7.085 1.1 6.365 1.1 6.365 0.5 5.805 0.5 5.805 1.58 5.645 1.58 5.645 1.8 5.525 1.8 5.525 1.46 5.685 1.46 5.685 0.38 6.485 0.38 6.485 0.98 6.965 0.98 6.965 0.48 6.845 0.48 6.845 0.36 7.085 0.36 ;
      POLYGON 6.245 1.1 6.045 1.1 6.045 1.92 6.11 1.92 6.11 2.04 5.125 2.04 5.125 1.58 4.865 1.58 4.865 1.42 4.745 1.42 4.745 1.3 4.985 1.3 4.985 1.46 5.245 1.46 5.245 1.92 5.925 1.92 5.925 0.98 6.125 0.98 6.125 0.62 6.245 0.62 ;
      POLYGON 5.325 0.48 5.225 0.48 5.225 0.96 4.505 0.96 4.505 0.56 3.995 0.56 3.995 0.765 4.115 0.765 4.115 1.825 3.685 1.825 3.685 1.965 3.565 1.965 3.565 1.705 3.995 1.705 3.995 0.885 3.875 0.885 3.875 0.44 4.625 0.44 4.625 0.84 5.105 0.84 5.105 0.48 5.085 0.48 5.085 0.36 5.325 0.36 ;
      POLYGON 3.315 0.505 3.195 0.505 3.195 1.125 2.595 1.125 2.595 0.525 2.235 0.525 2.235 1.86 2.115 1.86 2.115 0.64 1.815 0.64 1.815 0.4 1.935 0.4 1.935 0.405 2.715 0.405 2.715 1.005 3.075 1.005 3.075 0.385 3.315 0.385 ;
      POLYGON 2.625 2.25 1.555 2.25 1.555 2.13 2.505 2.13 2.505 1.965 2.355 1.965 2.355 0.645 2.475 0.645 2.475 1.845 2.625 1.845 ;
      POLYGON 1.435 1.48 1.315 1.48 1.315 1.68 0.595 1.68 0.595 1.86 0.475 1.86 0.475 1.74 0.135 1.74 0.135 0.4 0.255 0.4 0.255 1.56 1.195 1.56 1.195 1.36 1.435 1.36 ;
  END
END DLY3X1

MACRO OAI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X4 0 0 ;
  SIZE 11.02 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.96 1.06 6.36 1.18 ;
        RECT 4.945 1.23 5.205 1.38 ;
        RECT 4.96 1.06 5.205 1.38 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.295 1.06 9.56 1.3 ;
        RECT 9.295 1.06 9.555 1.38 ;
        RECT 8.1 1.06 9.56 1.18 ;
    END
  END C1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.31 1.06 2.83 1.18 ;
        RECT 1.465 1.06 1.725 1.38 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.03 1.175 7.18 1.435 ;
        RECT 4.18 1.5 7.15 1.62 ;
        RECT 7.03 1.175 7.15 1.62 ;
        RECT 5.325 1.3 5.565 1.62 ;
        RECT 4.18 1.22 4.3 1.62 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.61 1.5 9.88 1.62 ;
        RECT 9.76 1.22 9.88 1.62 ;
        RECT 8.72 1.3 8.96 1.62 ;
        RECT 7.61 1.175 7.76 1.62 ;
        RECT 7.46 1.28 7.76 1.4 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.432 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 1.5 3.41 1.62 ;
        RECT 3.26 1.175 3.41 1.62 ;
        RECT 1.97 1.3 2.21 1.62 ;
        RECT 0.57 1.28 0.69 1.62 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.7984 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.22 1.465 10.37 1.725 ;
        RECT 1.53 1.74 10.34 1.86 ;
        RECT 10.22 0.65 10.34 1.86 ;
        RECT 7.7 0.82 10.34 0.94 ;
        RECT 9.38 0.65 9.5 0.94 ;
        RECT 9.28 1.74 9.4 2.21 ;
        RECT 8.54 0.65 8.66 0.94 ;
        RECT 8 1.74 8.12 2.21 ;
        RECT 7.7 0.65 7.82 0.94 ;
        RECT 6.44 1.74 6.56 2.21 ;
        RECT 4.76 1.74 4.88 2.21 ;
        RECT 2.81 1.74 2.93 2.21 ;
        RECT 1.53 1.74 1.65 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 11.02 0.18 ;
        RECT 3.53 -0.18 3.65 0.7 ;
        RECT 2.69 -0.18 2.81 0.7 ;
        RECT 1.85 -0.18 1.97 0.7 ;
        RECT 1.01 -0.18 1.13 0.7 ;
        RECT 0.17 -0.18 0.29 0.7 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 11.02 2.79 ;
        RECT 9.86 1.98 10.1 2.15 ;
        RECT 9.86 1.98 9.98 2.79 ;
        RECT 8.58 1.98 8.82 2.15 ;
        RECT 8.58 1.98 8.7 2.79 ;
        RECT 7.22 1.98 7.46 2.15 ;
        RECT 7.22 1.98 7.34 2.79 ;
        RECT 5.605 1.98 5.845 2.15 ;
        RECT 5.605 1.98 5.725 2.79 ;
        RECT 3.86 1.98 4.1 2.15 ;
        RECT 3.86 1.98 3.98 2.79 ;
        RECT 2.11 1.98 2.35 2.15 ;
        RECT 2.11 1.98 2.23 2.79 ;
        RECT 0.89 1.74 1.01 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.76 0.7 10.64 0.7 10.64 0.53 9.92 0.53 9.92 0.7 9.8 0.7 9.8 0.53 9.08 0.53 9.08 0.7 8.96 0.7 8.96 0.53 8.24 0.53 8.24 0.7 8.12 0.7 8.12 0.53 7.4 0.53 7.4 0.7 7.28 0.7 7.28 0.53 6.56 0.53 6.56 0.7 6.44 0.7 6.44 0.53 5.72 0.53 5.72 0.7 5.6 0.7 5.6 0.53 4.88 0.53 4.88 0.7 4.76 0.7 4.76 0.53 4.04 0.53 4.04 0.7 3.92 0.7 3.92 0.41 10.76 0.41 ;
      POLYGON 6.98 0.94 0.59 0.94 0.59 0.65 0.71 0.65 0.71 0.82 1.43 0.82 1.43 0.65 1.55 0.65 1.55 0.82 2.27 0.82 2.27 0.65 2.39 0.65 2.39 0.82 3.11 0.82 3.11 0.65 3.23 0.65 3.23 0.82 4.34 0.82 4.34 0.65 4.46 0.65 4.46 0.82 5.18 0.82 5.18 0.65 5.3 0.65 5.3 0.82 6.02 0.82 6.02 0.65 6.14 0.65 6.14 0.82 6.86 0.82 6.86 0.65 6.98 0.65 ;
  END
END OAI222X4

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 1.45 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.216 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 1 0.49 1.24 ;
        RECT 0.07 1.025 0.49 1.145 ;
        RECT 0.07 0.885 0.22 1.145 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3456 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.885 0.8 1.145 ;
        RECT 0.65 0.68 0.77 2.01 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 1.45 0.18 ;
        RECT 1.07 -0.18 1.19 0.73 ;
        RECT 0.23 -0.18 0.35 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 1.45 2.79 ;
        RECT 1.07 1.36 1.19 2.79 ;
        RECT 0.23 1.36 0.35 2.79 ;
    END
  END VDD
END INVX2

MACRO TLATNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRXL 0 0 ;
  SIZE 7.83 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.945 1.25 2.065 1.49 ;
        RECT 1.755 1.52 2.015 1.67 ;
        RECT 1.895 1.37 2.015 1.67 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.98 1.12 5.175 1.495 ;
        RECT 4.98 1.12 5.12 1.5 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.67 1.255 6.91 1.375 ;
        RECT 6.19 1.175 6.79 1.295 ;
        RECT 6.19 0.885 6.475 1.295 ;
        RECT 6.355 0.375 6.475 1.295 ;
        RECT 5.425 0.375 6.475 0.495 ;
        RECT 6.16 0.885 6.475 1.145 ;
        RECT 4.775 0.64 5.545 0.76 ;
        RECT 5.425 0.375 5.545 0.76 ;
        RECT 4.775 0.36 4.895 0.76 ;
        RECT 3.065 0.36 4.895 0.48 ;
    END
  END RN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.03 1.175 7.335 1.415 ;
        RECT 7.03 1.175 7.18 1.435 ;
    END
  END GN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.68 0.255 1.58 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.365 1.585 1.485 1.83 ;
        RECT 1.365 0.65 1.485 0.89 ;
        RECT 1.23 1.465 1.445 1.725 ;
        RECT 1.325 0.77 1.445 1.725 ;
    END
  END QN
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 7.83 0.18 ;
        RECT 7.155 -0.18 7.275 0.795 ;
        RECT 5.185 -0.18 5.305 0.52 ;
        RECT 2.825 0.68 3.165 0.8 ;
        RECT 2.825 -0.18 2.945 0.8 ;
        RECT 1.785 -0.18 1.905 0.89 ;
        RECT 0.555 -0.18 0.675 0.92 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 7.83 2.79 ;
        RECT 7.03 1.655 7.15 2.79 ;
        RECT 6.19 1.655 6.31 2.79 ;
        RECT 5.065 1.62 5.185 2.79 ;
        RECT 3.525 1.89 3.645 2.79 ;
        RECT 2.685 2.23 2.805 2.79 ;
        RECT 1.845 2.23 1.965 2.79 ;
        RECT 0.615 1.98 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.695 0.935 7.575 0.935 7.575 1.655 7.57 1.655 7.57 1.775 7.45 1.775 7.45 1.535 7.455 1.535 7.455 1.055 6.595 1.055 6.595 0.935 7.455 0.935 7.455 0.815 7.575 0.815 7.575 0.555 7.695 0.555 ;
      POLYGON 6.73 1.775 6.61 1.775 6.61 1.655 6.43 1.655 6.43 1.535 5.92 1.535 5.92 1.24 5.545 1.24 5.545 1.12 5.92 1.12 5.92 0.615 6.235 0.615 6.235 0.735 6.04 0.735 6.04 1.415 6.55 1.415 6.55 1.535 6.73 1.535 ;
      POLYGON 5.785 1 5.425 1 5.425 1.5 5.605 1.5 5.605 1.74 5.485 1.74 5.485 1.62 5.305 1.62 5.305 1 4.845 1 4.845 1.12 4.185 1.12 4.185 1.2 3.945 1.2 3.945 1.08 4.065 1.08 4.065 1 4.725 1 4.725 0.88 5.665 0.88 5.665 0.62 5.785 0.62 ;
      POLYGON 4.605 0.88 3.825 0.88 3.825 1.32 4.445 1.32 4.445 1.74 4.325 1.74 4.325 1.44 2.425 1.44 2.425 1.32 3.705 1.32 3.705 0.76 4.485 0.76 4.485 0.62 4.605 0.62 ;
      POLYGON 4.085 1.68 3.965 1.68 3.965 1.77 2.985 1.77 2.985 1.65 3.845 1.65 3.845 1.56 4.085 1.56 ;
      POLYGON 3.585 1.2 3.465 1.2 3.465 1.13 2.305 1.13 2.305 1.59 2.325 1.59 2.325 1.83 2.205 1.83 2.205 1.71 2.185 1.71 2.185 1.13 1.805 1.13 1.805 1.17 1.565 1.17 1.565 1.01 2.425 1.01 2.425 0.65 2.545 0.65 2.545 1.01 3.465 1.01 3.465 0.96 3.585 0.96 ;
      POLYGON 1.095 1.58 0.975 1.58 0.975 1.2 0.375 1.2 0.375 1.08 0.975 1.08 0.975 0.68 1.095 0.68 ;
  END
END TLATNSRXL

MACRO MXI2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2XL 0 0 ;
  SIZE 2.32 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.15 1.265 0.27 1.595 ;
        RECT 0.07 1.1 0.22 1.435 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 1.44 1.4 1.85 ;
    END
  END B
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.55 1.2 1.74 1.44 ;
        RECT 1.52 1.465 1.67 1.725 ;
        RECT 1.55 1.2 1.67 1.725 ;
        RECT 0.87 1.2 1.74 1.32 ;
    END
  END S0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.192 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.39 0.72 0.96 0.84 ;
        RECT 0.78 1.89 0.9 2.13 ;
        RECT 0.39 1.89 0.9 2.01 ;
        RECT 0.39 0.72 0.51 2.01 ;
        RECT 0.36 0.885 0.51 1.145 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 2.32 0.18 ;
        RECT 1.37 0.72 1.61 0.84 ;
        RECT 1.37 -0.18 1.49 0.84 ;
        RECT 0.135 -0.18 0.255 0.38 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 2.32 2.79 ;
        RECT 1.42 1.97 1.54 2.79 ;
        RECT 0.14 1.97 0.26 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.98 1.68 1.96 1.68 1.96 2.09 1.84 2.09 1.84 1.56 1.86 1.56 1.86 1.08 0.75 1.08 0.75 1.44 1.04 1.44 1.04 1.77 0.92 1.77 0.92 1.56 0.63 1.56 0.63 0.96 1.08 0.96 1.08 0.6 0.68 0.6 0.68 0.5 0.56 0.5 0.56 0.38 0.8 0.38 0.8 0.48 1.25 0.48 1.25 0.96 1.85 0.96 1.85 0.66 1.97 0.66 1.97 0.78 1.98 0.78 ;
  END
END MXI2XL

MACRO OA22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X4 0 0 ;
  SIZE 4.35 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.94 1.175 1.235 1.295 ;
        RECT 1.115 1.055 1.235 1.295 ;
        RECT 0.94 1.175 1.09 1.435 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.01 0.51 1.465 ;
        RECT 0.38 1.01 0.5 1.495 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 1.03 0.82 1.435 ;
        RECT 0.7 1.02 0.82 1.435 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.81 1.465 1.96 1.725 ;
        RECT 1.81 1.34 1.93 1.725 ;
        RECT 1.6 1.34 1.93 1.46 ;
        RECT 1.6 1.22 1.72 1.46 ;
    END
  END B0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 1.175 3.7 1.435 ;
        RECT 2.685 0.74 3.585 0.86 ;
        RECT 3.465 0.62 3.585 0.86 ;
        RECT 2.08 1.32 3.525 1.44 ;
        RECT 3.405 0.74 3.525 1.44 ;
        RECT 2.92 1.32 3.04 2.21 ;
        RECT 2.565 0.69 2.805 0.81 ;
        RECT 2.08 1.32 2.2 2.21 ;
    END
  END Y
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 4.35 0.18 ;
        RECT 3.885 -0.18 4.005 0.68 ;
        RECT 2.985 0.5 3.225 0.62 ;
        RECT 2.985 -0.18 3.105 0.62 ;
        RECT 2.205 -0.18 2.325 0.68 ;
        RECT 0.555 -0.18 0.675 0.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 4.35 2.79 ;
        RECT 3.34 1.56 3.46 2.79 ;
        RECT 2.5 1.56 2.62 2.79 ;
        RECT 1.66 1.845 1.78 2.79 ;
        RECT 0.22 1.615 0.34 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 3.285 1.15 3.045 1.15 3.045 1.1 2.54 1.1 2.54 1.13 2.3 1.13 2.3 1.1 1.48 1.1 1.48 1.675 1.095 1.675 1.095 2.21 0.975 2.21 0.975 1.555 1.36 1.555 1.36 0.72 1.395 0.72 1.395 0.6 1.515 0.6 1.515 0.84 1.48 0.84 1.48 0.98 3.165 0.98 3.165 1.03 3.285 1.03 ;
      POLYGON 1.935 0.65 1.815 0.65 1.815 0.48 1.095 0.48 1.095 0.89 0.135 0.89 0.135 0.6 0.255 0.6 0.255 0.77 0.975 0.77 0.975 0.36 1.935 0.36 ;
  END
END OA22X4

MACRO DFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX8 0 0 ;
  SIZE 9.57 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.53 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.655 0.68 2.775 2.13 ;
        RECT 0.07 1.025 2.775 1.145 ;
        RECT 1.815 0.68 1.935 2.13 ;
        RECT 0.975 0.68 1.095 2.125 ;
        RECT 0.135 0.68 0.255 2.125 ;
        RECT 0.07 0.885 0.255 1.145 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.086 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.77 1.06 8.92 1.435 ;
        RECT 8.725 1.04 8.845 1.425 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.04 1.04 9.215 1.45 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 9.57 0.18 ;
        RECT 8.885 -0.18 9.005 0.68 ;
        RECT 7.325 0.4 7.565 0.52 ;
        RECT 7.325 -0.18 7.445 0.52 ;
        RECT 5.485 0.5 5.725 0.62 ;
        RECT 5.485 -0.18 5.605 0.62 ;
        RECT 3.915 -0.18 4.035 0.73 ;
        RECT 3.075 -0.18 3.195 0.73 ;
        RECT 2.235 -0.18 2.355 0.67 ;
        RECT 1.395 -0.18 1.515 0.67 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 9.57 2.79 ;
        RECT 8.585 1.81 8.825 1.93 ;
        RECT 8.585 1.81 8.705 2.79 ;
        RECT 7.245 2.08 7.485 2.2 ;
        RECT 7.245 2.08 7.365 2.79 ;
        RECT 5.265 2.26 5.505 2.79 ;
        RECT 3.915 2.02 4.155 2.14 ;
        RECT 3.915 2.02 4.035 2.79 ;
        RECT 3.075 1.48 3.195 2.79 ;
        RECT 2.235 1.385 2.355 2.79 ;
        RECT 1.395 1.385 1.515 2.79 ;
        RECT 0.555 1.385 0.675 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 9.425 0.8 9.245 0.8 9.245 0.92 8.525 0.92 8.525 1.57 9.325 1.57 9.325 1.81 9.205 1.81 9.205 1.69 8.465 1.69 8.465 2.23 8.045 2.23 8.045 2.25 7.805 2.25 7.805 2.23 7.645 2.23 7.645 1.96 6.705 1.96 6.705 2.23 5.625 2.23 5.625 2.14 4.945 2.14 4.945 2.02 5.745 2.02 5.745 2.11 6.585 2.11 6.585 1.24 6.745 1.24 6.745 1.12 6.865 1.12 6.865 1.36 6.705 1.36 6.705 1.84 7.765 1.84 7.765 2.11 8.345 2.11 8.345 1.57 8.405 1.57 8.405 0.8 9.125 0.8 9.125 0.68 9.305 0.68 9.305 0.44 9.425 0.44 ;
      POLYGON 8.305 0.68 8.285 0.68 8.285 1.36 8.125 1.36 8.125 1.99 8.005 1.99 8.005 1.36 7.345 1.36 7.345 1.31 7.225 1.31 7.225 1.19 7.465 1.19 7.465 1.24 8.165 1.24 8.165 0.56 8.185 0.56 8.185 0.44 8.305 0.44 ;
      POLYGON 8.045 1.12 7.925 1.12 7.925 0.76 7.085 0.76 7.085 0.48 6.605 0.48 6.605 1.12 6.405 1.12 6.405 0.88 6.485 0.88 6.485 0.48 6.005 0.48 6.005 0.86 5.985 0.86 5.985 1.53 5.025 1.53 5.025 1.65 4.785 1.65 4.785 1.53 4.905 1.53 4.905 1.41 5.865 1.41 5.865 0.86 5.065 0.86 5.065 0.54 5.185 0.54 5.185 0.74 5.885 0.74 5.885 0.36 7.205 0.36 7.205 0.64 8.045 0.64 ;
      POLYGON 7.785 1.07 7.105 1.07 7.105 1.6 6.945 1.6 6.945 1.72 6.825 1.72 6.825 1.48 6.985 1.48 6.985 1 6.725 1 6.725 0.6 6.965 0.6 6.965 0.88 7.105 0.88 7.105 0.95 7.785 0.95 ;
      POLYGON 6.365 0.72 6.245 0.72 6.245 1.99 6.125 1.99 6.125 1.9 4.155 1.9 4.155 1.34 4.035 1.34 4.035 1.22 4.275 1.22 4.275 1.78 6.125 1.78 6.125 0.6 6.365 0.6 ;
      POLYGON 5.725 1.1 4.515 1.1 4.515 1.54 4.635 1.54 4.635 1.66 4.395 1.66 4.395 1.1 3.615 1.1 3.615 2.13 3.495 2.13 3.495 1.1 3.055 1.1 3.055 1.24 2.935 1.24 2.935 0.98 3.495 0.98 3.495 0.68 3.615 0.68 3.615 0.98 4.335 0.98 4.335 0.68 4.455 0.68 4.455 0.8 4.515 0.8 4.515 0.98 5.725 0.98 ;
  END
END DFFHQX8

MACRO EDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX4 0 0 ;
  SIZE 10.15 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 1.06 0.51 1.515 ;
        RECT 0.36 1.03 0.48 1.515 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.108 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.06 1.03 9.24 1.45 ;
        RECT 9.12 1.01 9.24 1.45 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.168 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.585 1.23 9.845 1.38 ;
        RECT 9.5 1.14 9.705 1.26 ;
        RECT 9.5 0.77 9.62 1.26 ;
        RECT 8.82 0.77 9.62 0.89 ;
        RECT 8.7 0.98 8.94 1.1 ;
        RECT 8.82 0.36 8.94 1.1 ;
        RECT 8.22 0.36 8.94 0.48 ;
        RECT 8.22 0.36 8.34 1.08 ;
        RECT 8.18 0.96 8.3 1.44 ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.7944 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.145 0.65 6.385 0.77 ;
        RECT 6.025 1.58 6.265 1.71 ;
        RECT 5.065 0.94 6.265 1.06 ;
        RECT 6.145 0.65 6.265 1.06 ;
        RECT 5.065 1.58 6.265 1.7 ;
        RECT 5.125 1.47 5.245 1.71 ;
        RECT 5.065 0.65 5.185 1.7 ;
        RECT 4.945 1.52 5.245 1.67 ;
        RECT 4.945 0.65 5.185 0.77 ;
    END
  END Q
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 10.15 0.18 ;
        RECT 9.26 -0.18 9.38 0.65 ;
        RECT 7.645 -0.18 7.765 0.45 ;
        RECT 6.745 -0.18 6.865 0.64 ;
        RECT 5.545 0.46 5.785 0.58 ;
        RECT 5.665 -0.18 5.785 0.58 ;
        RECT 4.465 -0.18 4.585 0.68 ;
        RECT 2.625 0.43 2.865 0.55 ;
        RECT 2.745 -0.18 2.865 0.55 ;
        RECT 0.555 -0.18 0.675 0.67 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 10.15 2.79 ;
        RECT 9.26 1.81 9.38 2.79 ;
        RECT 7.525 2.16 7.645 2.79 ;
        RECT 6.565 2.07 6.685 2.79 ;
        RECT 5.545 2.07 5.785 2.19 ;
        RECT 5.545 2.07 5.665 2.79 ;
        RECT 4.585 2.07 4.825 2.19 ;
        RECT 4.585 2.07 4.705 2.79 ;
        RECT 2.745 1.75 2.865 2.79 ;
        RECT 0.615 2.155 0.735 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 10.085 1.69 9.86 1.69 9.86 1.81 9.74 1.81 9.74 1.69 8.82 1.69 8.82 1.42 8.7 1.42 8.7 1.3 8.94 1.3 8.94 1.57 9.965 1.57 9.965 1.02 9.74 1.02 9.74 0.6 9.86 0.6 9.86 0.9 10.085 0.9 ;
      POLYGON 8.7 0.86 8.58 0.86 8.58 2.21 8.46 2.21 8.46 2.04 7.665 2.04 7.665 1.95 4.215 1.95 4.215 2.23 3.035 2.23 3.035 1.63 2.625 1.63 2.625 2.23 1.445 2.23 1.445 1.59 1.345 1.59 1.345 0.72 1.305 0.72 1.305 0.6 1.545 0.6 1.545 0.72 1.465 0.72 1.465 1.47 1.565 1.47 1.565 2.11 2.505 2.11 2.505 1.51 3.155 1.51 3.155 2.11 4.095 2.11 4.095 1.83 7.785 1.83 7.785 1.92 8.46 1.92 8.46 0.74 8.58 0.74 8.58 0.6 8.7 0.6 ;
      POLYGON 8.16 1.8 8.04 1.8 8.04 1.68 7.94 1.68 7.94 1.56 7.165 1.56 7.165 1.71 7.045 1.71 7.045 1.46 5.885 1.46 5.885 1.21 6.125 1.21 6.125 1.34 7.405 1.34 7.405 0.78 7.165 0.78 7.165 0.5 7.285 0.5 7.285 0.66 7.525 0.66 7.525 0.72 7.98 0.72 7.98 0.6 8.1 0.6 8.1 0.84 7.525 0.84 7.525 1.44 8.06 1.44 8.06 1.56 8.16 1.56 ;
      POLYGON 7.285 1.02 6.945 1.02 6.945 1.22 6.705 1.22 6.705 1.1 6.825 1.1 6.825 0.88 6.505 0.88 6.505 0.53 6.025 0.53 6.025 0.82 5.305 0.82 5.305 0.53 4.825 0.53 4.825 0.92 4.465 0.92 4.465 1.61 4.125 1.61 4.125 1.71 3.885 1.71 3.885 1.53 4.005 1.53 4.005 1.49 4.345 1.49 4.345 0.92 3.825 0.92 3.825 0.54 3.945 0.54 3.945 0.8 4.705 0.8 4.705 0.41 5.425 0.41 5.425 0.7 5.905 0.7 5.905 0.41 6.625 0.41 6.625 0.76 6.945 0.76 6.945 0.9 7.285 0.9 ;
      POLYGON 4.225 1.37 4.105 1.37 4.105 1.25 3.585 1.25 3.585 1.12 3.565 1.12 3.565 0.88 3.585 0.88 3.585 0.48 3.105 0.48 3.105 0.79 2.385 0.79 2.385 1.12 2.145 1.12 2.145 0.88 2.265 0.88 2.265 0.48 1.785 0.48 1.785 0.96 1.705 0.96 1.705 1.35 1.585 1.35 1.585 0.84 1.665 0.84 1.665 0.48 1.185 0.48 1.185 1.635 1.175 1.635 1.175 1.755 1.055 1.755 1.055 1.515 1.065 1.515 1.065 0.67 0.975 0.67 0.975 0.36 2.505 0.36 2.505 0.67 2.985 0.67 2.985 0.36 3.705 0.36 3.705 1.13 4.225 1.13 ;
      POLYGON 3.465 0.72 3.445 0.72 3.445 1.39 3.395 1.39 3.395 1.99 3.275 1.99 3.275 1.39 2.745 1.39 2.745 1.15 2.865 1.15 2.865 1.27 3.325 1.27 3.325 0.72 3.225 0.72 3.225 0.6 3.465 0.6 ;
      POLYGON 3.205 1.15 3.085 1.15 3.085 1.03 2.625 1.03 2.625 1.36 2.025 1.36 2.025 1.99 1.905 1.99 1.905 0.6 2.145 0.6 2.145 0.72 2.025 0.72 2.025 1.24 2.505 1.24 2.505 0.91 3.205 0.91 ;
      POLYGON 0.945 0.95 0.705 0.95 0.705 0.91 0.24 0.91 0.24 1.635 0.255 1.635 0.255 1.875 0.135 1.875 0.135 1.755 0.12 1.755 0.12 0.67 0.135 0.67 0.135 0.43 0.255 0.43 0.255 0.79 0.945 0.79 ;
  END
END EDFFHQX4

MACRO TLATNCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX4 0 0 ;
  SIZE 6.38 BY 2.61 ;
  SYMMETRY X Y ;
  SITE gsclib090site ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.885 0.835 1.185 ;
        RECT 0.61 0.955 0.77 1.24 ;
    END
  END CK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.525 1.22 5.785 1.44 ;
        RECT 5.525 1.22 5.645 1.57 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.6912 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 1.4 2.275 1.58 ;
        RECT 2.015 0.74 2.255 0.86 ;
        RECT 1.235 0.79 2.135 0.91 ;
        RECT 1.23 1.3 2.155 1.42 ;
        RECT 1.23 1.175 1.38 1.435 ;
        RECT 1.235 0.67 1.355 1.46 ;
        RECT 1.135 1.34 1.255 1.58 ;
    END
  END ECK
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.18 6.38 0.18 ;
        RECT 5.525 0.5 5.765 0.62 ;
        RECT 5.645 -0.18 5.765 0.62 ;
        RECT 4.005 0.62 4.125 0.86 ;
        RECT 3.965 -0.18 4.085 0.74 ;
        RECT 2.495 -0.18 2.615 0.73 ;
        RECT 1.595 0.55 1.835 0.67 ;
        RECT 1.595 -0.18 1.715 0.67 ;
        RECT 0.815 -0.18 0.935 0.73 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 2.43 6.38 2.79 ;
        RECT 5.605 1.69 5.725 2.79 ;
        RECT 4.205 2.1 4.445 2.22 ;
        RECT 4.205 2.1 4.325 2.79 ;
        RECT 3.305 2.12 3.425 2.79 ;
        RECT 2.575 2.12 2.695 2.79 ;
        RECT 1.555 1.94 1.795 2.06 ;
        RECT 1.555 1.94 1.675 2.79 ;
        RECT 0.655 1.94 0.775 2.79 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 6.265 1.75 5.965 1.75 5.965 1.63 6.145 1.63 6.145 0.86 5.285 0.86 5.285 0.48 4.205 0.48 4.205 0.36 5.405 0.36 5.405 0.74 6.065 0.74 6.065 0.62 6.185 0.62 6.185 0.74 6.265 0.74 ;
      POLYGON 6.025 1.22 5.905 1.22 5.905 1.1 5.405 1.1 5.405 1.71 5.145 1.71 5.145 1.75 4.905 1.75 4.905 1.63 5.025 1.63 5.025 1.59 5.285 1.59 5.285 1.1 4.765 1.1 4.765 0.62 4.885 0.62 4.885 0.98 6.025 0.98 ;
      POLYGON 5.165 1.47 5.045 1.47 5.045 1.35 3.235 1.35 3.235 1.52 2.995 1.52 2.995 1.4 3.115 1.4 3.115 0.92 2.975 0.92 2.975 0.68 3.095 0.68 3.095 0.8 3.235 0.8 3.235 1.23 4.505 1.23 4.505 0.96 4.625 0.96 4.625 1.23 5.165 1.23 ;
      POLYGON 4.945 2.25 4.825 2.25 4.825 1.99 4.565 1.99 4.565 1.98 3.89 1.98 3.89 2 2.445 2 2.445 1.82 0.175 1.82 0.175 1.46 0.335 1.46 0.335 0.68 0.455 0.68 0.455 1.58 0.295 1.58 0.295 1.7 2.565 1.7 2.565 1.88 3.77 1.88 3.77 1.86 4.685 1.86 4.685 1.87 4.945 1.87 ;
      POLYGON 3.965 1.74 3.58 1.74 3.58 1.76 2.735 1.76 2.735 1.18 1.895 1.18 1.895 1.06 2.735 1.06 2.735 0.44 3.485 0.44 3.485 0.73 3.365 0.73 3.365 0.56 2.855 0.56 2.855 1.64 3.46 1.64 3.46 1.62 3.965 1.62 ;
  END
END TLATNCAX4

END LIBRARY
