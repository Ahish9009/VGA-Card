module pixel_itr(
    input wire clk,
    input wire pix_clk,
    input wire rst,
    output wire [9:0] pix_x,
    output wire [9:0] pix_y,
    output wire h_sync,
    output wire v_sync,
    output wire draw_active,
    output wire screen_end,
    output wire draw_end
    );
	 
	// FOR 800 X 600
    // parameter h_sync_strt = 56;          
    // parameter h_sync_end  = 56 + 120;         
    // parameter v_sync_strt = 600 + 37;        
    // parameter v_sync_end  = 600 + 37 + 6;   
    // parameter h_draw_min  = 56 + 120 + 64;   
    // parameter v_draw_max  = 600 - 1;            
    // parameter h_max = 1040;           
    // parameter v_max = 666 - 1;
	 
	// FOR 640 X 480
    parameter h_sync_strt = 16;          
    parameter h_sync_end  = 16 + 96;         
    parameter v_sync_strt = 480 + 10;        
    parameter v_sync_end  = 480 + 10 + 2;   
    parameter h_draw_min  = 16 + 96 + 48;   
    parameter v_draw_max  = 480 - 1;            
    parameter h_max = 800;           
    parameter v_max = 525 - 1;

    reg [9:0] h_pos=0;
	 reg [9:0] v_pos=0; 
	
    // --------------- SYNC SIGNALS BLOCK ---------------
    assign h_sync = (h_pos >= h_sync_strt && h_pos < h_sync_end) ? 0 : 1;
    assign v_sync = (v_pos >= v_sync_strt && v_pos < v_sync_end) ? 0 : 1;
    // --------------------------------------------------
		
	// -------------- PIXEL POSITION BLOCK --------------
    // assign pix_x = (h_pos >= h_draw_min) ? h_pos : 0;        
    assign pix_x = (h_pos >= h_draw_min) ? h_pos - h_draw_min : 0;        
	 assign pix_y = (v_pos <= v_draw_max) ? v_pos : v_draw_max;        
    // --------------------------------------------------

    // -------- BLANKING / DRAWING PERIOD BLOCK ---------
    assign draw_active = (h_pos < h_draw_min | v_pos > v_draw_max) ? 0 : 1;
    // --------------------------------------------------

    // ----------------- LIMITS BLOCK -------------------
    assign screen_end = (h_pos == h_max & v_pos == v_max);
    assign draw_end = (h_pos == h_max & v_pos == v_draw_max);
    // --------------------------------------------------
    
    // ------------------ MAIN BLOCK --------------------
    always @ (posedge clk) begin
        if (rst) begin
            h_pos <= 0; 
            v_pos <= 0;
        end

        if(pix_clk) begin
            if (h_pos < h_max) begin
                h_pos <= h_pos + 1; 
            end
            else begin
                h_pos <= 0;
                v_pos <= v_pos + 1;
            end

            if (v_pos == v_max) begin
                    v_pos <= 0;
            end
        end
    end
    // --------------------------------------------------

endmodule

//////////////////////////////////////////////////////////////////////////////////

module screen_design(
	input clk,
	input rst,
	output h_sync,
	output v_sync,
	output r_out,
	output g_out,
	output b_out
);

//---------------GENERATING PIXEL CLOCK----------------------
reg count = 0, pix_clk = 0;

always @(posedge clk) begin
	
	if (rst == 1) begin
		count <= 0;
		pix_clk <= 0;
	end 
	if (count == 1) begin
		pix_clk <= 1;
		count <= 0;
	end 
	else begin
		pix_clk <= 0;
		count <= count + 1;

	end
end

//-----------------------------------------------------------

//-------------GETTING CURRENT PIXEL COORDINATES-------------
wire [9:0] pix_x;
wire [9:0] pix_y;

pixel_itr show(
	.clk(clk),
   .pix_clk(pix_clk),
	.rst(rst),
	.pix_x(pix_x),
	.pix_y(pix_y),
	.h_sync(h_sync),
	.v_sync(v_sync)
);
//-----------------------------------------------------------

//----------GENERATING WINDOWS LOGO(4 SQUARES)---------------



//---------RED---------


assign r_out =  (pix_x >= 404 & pix_x <=405 & pix_y >= 111 & pix_y <=111 ) | (pix_x >= 409 & pix_x <=410 & pix_y >= 111 & pix_y <=111 ) | (pix_x >= 393 & pix_x <=400 & pix_y >= 112 & pix_y <=112 ) | (pix_x >= 403 & pix_x <=413 & pix_y >= 112 & pix_y <=112 ) | (pix_x >= 391 & pix_x <=426 & pix_y >= 113 & pix_y <=113 ) | (pix_x >= 387 & pix_x <=427 & pix_y >= 114 & pix_y <=114 ) | (pix_x >= 384 & pix_x <=428 & pix_y >= 115 & pix_y <=115 ) | (pix_x >= 382 & pix_x <=428 & pix_y >= 116 & pix_y <=116 ) | (pix_x >= 380 & pix_x <=429 & pix_y >= 117 & pix_y <=117 ) | (pix_x >= 376 & pix_x <=430 & pix_y >= 118 & pix_y <=118 ) | (pix_x >= 375 & pix_x <=431 & pix_y >= 119 & pix_y <=119 ) | (pix_x >= 377 & pix_x <=431 & pix_y >= 120 & pix_y <=120 ) | (pix_x >= 377 & pix_x <=431 & pix_y >= 121 & pix_y <=121 ) | (pix_x >= 435 & pix_x <=436 & pix_y >= 121 & pix_y <=121 ) | (pix_x >= 375 & pix_x <=437 & pix_y >= 122 & pix_y <=122 ) | (pix_x >= 375 & pix_x <=438 & pix_y >= 123 & pix_y <=123 ) | (pix_x >= 375 & pix_x <=438 & pix_y >= 124 & pix_y <=124 ) | (pix_x >= 375 & pix_x <=437 & pix_y >= 125 & pix_y <=125 ) | (pix_x >= 377 & pix_x <=437 & pix_y >= 126 & pix_y <=126 ) | (pix_x >= 377 & pix_x <=438 & pix_y >= 127 & pix_y <=127 ) | (pix_x >= 376 & pix_x <=438 & pix_y >= 128 & pix_y <=127 ) | (pix_x >= 378 & pix_x <=438 & pix_y >= 128 & pix_y <=128 ) | (pix_x >= 376 & pix_x <=438 & pix_y >= 129 & pix_y <=128 ) | (pix_x >= 378 & pix_x <=439 & pix_y >= 129 & pix_y <=129 ) | (pix_x >= 376 & pix_x <=439 & pix_y >= 130 & pix_y <=129 ) | (pix_x >= 378 & pix_x <=441 & pix_y >= 130 & pix_y <=130 ) | (pix_x >= 376 & pix_x <=442 & pix_y >= 131 & pix_y <=131 ) | (pix_x >= 376 & pix_x <=443 & pix_y >= 132 & pix_y <=132 ) | (pix_x >= 377 & pix_x <=444 & pix_y >= 133 & pix_y <=133 ) | (pix_x >= 377 & pix_x <=446 & pix_y >= 134 & pix_y <=134 ) | (pix_x >= 377 & pix_x <=446 & pix_y >= 135 & pix_y <=135 ) | (pix_x >= 375 & pix_x <=448 & pix_y >= 136 & pix_y <=136 ) | (pix_x >= 375 & pix_x <=448 & pix_y >= 137 & pix_y <=137 ) | (pix_x >= 374 & pix_x <=448 & pix_y >= 138 & pix_y <=138 ) | (pix_x >= 374 & pix_x <=449 & pix_y >= 139 & pix_y <=139 ) | (pix_x >= 374 & pix_x <=449 & pix_y >= 140 & pix_y <=140 ) | (pix_x >= 374 & pix_x <=449 & pix_y >= 141 & pix_y <=141 ) | (pix_x >= 375 & pix_x <=450 & pix_y >= 142 & pix_y <=142 ) | (pix_x >= 375 & pix_x <=450 & pix_y >= 143 & pix_y <=143 ) | (pix_x >= 373 & pix_x <=451 & pix_y >= 144 & pix_y <=144 ) | (pix_x >= 374 & pix_x <=451 & pix_y >= 145 & pix_y <=145 ) | (pix_x >= 374 & pix_x <=452 & pix_y >= 146 & pix_y <=146 ) | (pix_x >= 373 & pix_x <=452 & pix_y >= 147 & pix_y <=147 ) | (pix_x >= 371 & pix_x <=453 & pix_y >= 148 & pix_y <=148 ) | (pix_x >= 371 & pix_x <=454 & pix_y >= 149 & pix_y <=149 ) | (pix_x >= 369 & pix_x <=454 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 369 & pix_x <=454 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 367 & pix_x <=403 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 411 & pix_x <=455 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 366 & pix_x <=400 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 408 & pix_x <=456 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 364 & pix_x <=397 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 406 & pix_x <=456 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 363 & pix_x <=395 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 404 & pix_x <=456 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 361 & pix_x <=387 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 403 & pix_x <=457 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 361 & pix_x <=386 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 403 & pix_x <=457 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 361 & pix_x <=384 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 404 & pix_x <=458 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 360 & pix_x <=384 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 400 & pix_x <=384 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 404 & pix_x <=416 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 419 & pix_x <=416 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 433 & pix_x <=458 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 358 & pix_x <=384 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 401 & pix_x <=420 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 433 & pix_x <=459 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 357 & pix_x <=384 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 400 & pix_x <=424 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 438 & pix_x <=459 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 356 & pix_x <=384 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 399 & pix_x <=422 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 355 & pix_x <=384 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 398 & pix_x <=420 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 353 & pix_x <=384 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 398 & pix_x <=422 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 353 & pix_x <=382 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 398 & pix_x <=422 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 353 & pix_x <=380 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 398 & pix_x <=424 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 353 & pix_x <=378 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 393 & pix_x <=394 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 398 & pix_x <=430 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 351 & pix_x <=376 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 391 & pix_x <=392 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 396 & pix_x <=392 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 410 & pix_x <=435 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 350 & pix_x <=372 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 410 & pix_x <=440 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 350 & pix_x <=368 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 436 & pix_x <=442 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 349 & pix_x <=368 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 348 & pix_x <=360 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 347 & pix_x <=351 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 445 & pix_x <=458 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 411 & pix_x <=416 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 447 & pix_x <=456 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 412 & pix_x <=433 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 448 & pix_x <=456 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 414 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 444 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 450 & pix_x <=456 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 414 & pix_x <=432 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 451 & pix_x <=455 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 404 & pix_x <=405 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 419 & pix_x <=416 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 453 & pix_x <=455 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 423 & pix_x <=433 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 453 & pix_x <=454 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 278 & pix_x <=280 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 363 & pix_x <=384 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 423 & pix_x <=431 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 433 & pix_x <=431 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 278 & pix_x <=281 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 356 & pix_x <=383 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 385 & pix_x <=383 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 415 & pix_x <=416 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 422 & pix_x <=431 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 433 & pix_x <=431 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 279 & pix_x <=282 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 350 & pix_x <=387 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 421 & pix_x <=433 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 443 & pix_x <=449 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 456 & pix_x <=458 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 279 & pix_x <=283 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 348 & pix_x <=387 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 423 & pix_x <=433 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 456 & pix_x <=458 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 281 & pix_x <=284 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 347 & pix_x <=387 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 407 & pix_x <=408 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 281 & pix_x <=284 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 347 & pix_x <=387 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 465 & pix_x <=468 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 281 & pix_x <=284 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 348 & pix_x <=387 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 463 & pix_x <=469 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 349 & pix_x <=388 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 455 & pix_x <=458 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 463 & pix_x <=464 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 350 & pix_x <=389 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 400 & pix_x <=408 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 351 & pix_x <=392 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 399 & pix_x <=408 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 352 & pix_x <=394 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 398 & pix_x <=408 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 422 & pix_x <=418 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 353 & pix_x <=408 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 422 & pix_x <=418 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 454 & pix_x <=455 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 462 & pix_x <=467 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 349 & pix_x <=409 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 421 & pix_x <=422 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 425 & pix_x <=434 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 442 & pix_x <=446 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 454 & pix_x <=456 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 258 & pix_x <=466 & pix_y >= 193 & pix_y <=192 ) | (pix_x >= 349 & pix_x <=351 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 415 & pix_x <=422 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 425 & pix_x <=436 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 442 & pix_x <=446 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 454 & pix_x <=457 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 415 & pix_x <=423 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 425 & pix_x <=437 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 442 & pix_x <=446 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 454 & pix_x <=459 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 415 & pix_x <=438 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 442 & pix_x <=446 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 453 & pix_x <=460 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 354 & pix_x <=409 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 442 & pix_x <=445 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 355 & pix_x <=409 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 445 & pix_x <=446 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 355 & pix_x <=409 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 445 & pix_x <=446 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 448 & pix_x <=449 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 355 & pix_x <=409 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 441 & pix_x <=449 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 356 & pix_x <=409 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 441 & pix_x <=448 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 452 & pix_x <=467 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 355 & pix_x <=409 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 441 & pix_x <=447 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 452 & pix_x <=467 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 355 & pix_x <=409 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 441 & pix_x <=447 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 452 & pix_x <=468 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 256 & pix_x <=260 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 354 & pix_x <=409 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 441 & pix_x <=446 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 452 & pix_x <=469 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 441 & pix_x <=446 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 451 & pix_x <=470 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 441 & pix_x <=446 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 451 & pix_x <=471 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 441 & pix_x <=445 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 451 & pix_x <=472 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 416 & pix_x <=445 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 451 & pix_x <=472 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 450 & pix_x <=474 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 450 & pix_x <=474 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 353 & pix_x <=409 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 441 & pix_x <=443 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 450 & pix_x <=476 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 353 & pix_x <=410 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 441 & pix_x <=443 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 449 & pix_x <=476 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 256 & pix_x <=259 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 353 & pix_x <=410 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 417 & pix_x <=443 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 449 & pix_x <=477 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 355 & pix_x <=360 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 362 & pix_x <=411 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 418 & pix_x <=440 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 449 & pix_x <=478 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 257 & pix_x <=259 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 356 & pix_x <=360 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 363 & pix_x <=411 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 419 & pix_x <=440 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 449 & pix_x <=480 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 267 & pix_x <=270 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 356 & pix_x <=360 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 364 & pix_x <=412 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 420 & pix_x <=440 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 449 & pix_x <=480 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 267 & pix_x <=271 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 361 & pix_x <=413 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 421 & pix_x <=439 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 447 & pix_x <=481 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 257 & pix_x <=260 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 268 & pix_x <=271 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 361 & pix_x <=414 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 422 & pix_x <=439 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 446 & pix_x <=481 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 258 & pix_x <=261 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 268 & pix_x <=271 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 361 & pix_x <=416 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 424 & pix_x <=439 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 444 & pix_x <=482 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 258 & pix_x <=261 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 268 & pix_x <=272 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 362 & pix_x <=418 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 426 & pix_x <=439 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 449 & pix_x <=483 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 259 & pix_x <=262 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 269 & pix_x <=272 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 362 & pix_x <=420 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 428 & pix_x <=442 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 448 & pix_x <=483 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 259 & pix_x <=262 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 269 & pix_x <=272 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 363 & pix_x <=422 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 431 & pix_x <=440 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 447 & pix_x <=484 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 260 & pix_x <=263 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 270 & pix_x <=273 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 363 & pix_x <=425 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 447 & pix_x <=484 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 260 & pix_x <=263 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 270 & pix_x <=274 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 363 & pix_x <=368 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 370 & pix_x <=429 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 449 & pix_x <=485 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 261 & pix_x <=264 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 271 & pix_x <=275 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 369 & pix_x <=432 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 447 & pix_x <=485 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 261 & pix_x <=264 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 271 & pix_x <=276 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 369 & pix_x <=431 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 447 & pix_x <=485 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 262 & pix_x <=266 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 272 & pix_x <=277 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 369 & pix_x <=429 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 449 & pix_x <=485 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 262 & pix_x <=266 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 273 & pix_x <=278 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 369 & pix_x <=428 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 433 & pix_x <=436 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 449 & pix_x <=486 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 263 & pix_x <=267 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 274 & pix_x <=280 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 369 & pix_x <=437 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 450 & pix_x <=486 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 263 & pix_x <=269 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 273 & pix_x <=285 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 370 & pix_x <=437 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 451 & pix_x <=485 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 263 & pix_x <=271 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 273 & pix_x <=288 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 370 & pix_x <=436 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 451 & pix_x <=485 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 264 & pix_x <=271 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 273 & pix_x <=278 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 282 & pix_x <=288 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 370 & pix_x <=436 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 451 & pix_x <=485 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 265 & pix_x <=274 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 282 & pix_x <=290 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 370 & pix_x <=436 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 452 & pix_x <=472 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 474 & pix_x <=485 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 265 & pix_x <=274 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 283 & pix_x <=292 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 370 & pix_x <=436 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 454 & pix_x <=463 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 474 & pix_x <=485 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 265 & pix_x <=275 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 285 & pix_x <=294 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 370 & pix_x <=436 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 455 & pix_x <=461 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 475 & pix_x <=484 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 267 & pix_x <=276 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 280 & pix_x <=276 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 286 & pix_x <=294 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 371 & pix_x <=437 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 454 & pix_x <=459 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 475 & pix_x <=484 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 267 & pix_x <=281 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 286 & pix_x <=296 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 371 & pix_x <=437 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 453 & pix_x <=457 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 476 & pix_x <=484 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 268 & pix_x <=296 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 371 & pix_x <=437 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 453 & pix_x <=456 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 476 & pix_x <=483 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 269 & pix_x <=296 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 371 & pix_x <=437 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 453 & pix_x <=455 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 477 & pix_x <=483 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 270 & pix_x <=296 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 371 & pix_x <=437 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 477 & pix_x <=482 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 270 & pix_x <=296 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 373 & pix_x <=438 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 452 & pix_x <=458 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 477 & pix_x <=481 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 271 & pix_x <=296 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 373 & pix_x <=438 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 451 & pix_x <=462 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 478 & pix_x <=462 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 272 & pix_x <=296 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 374 & pix_x <=439 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 451 & pix_x <=462 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 273 & pix_x <=296 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 377 & pix_x <=440 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 452 & pix_x <=462 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 274 & pix_x <=297 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 377 & pix_x <=444 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 451 & pix_x <=463 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 275 & pix_x <=298 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 377 & pix_x <=464 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 276 & pix_x <=298 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 375 & pix_x <=465 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 276 & pix_x <=298 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 375 & pix_x <=468 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 278 & pix_x <=300 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 375 & pix_x <=468 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 278 & pix_x <=301 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 375 & pix_x <=467 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 279 & pix_x <=301 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 374 & pix_x <=467 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 281 & pix_x <=301 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 374 & pix_x <=467 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 281 & pix_x <=300 & pix_y >= 252 & pix_y <=252 ) | (pix_x >= 374 & pix_x <=467 & pix_y >= 252 & pix_y <=252 ) | (pix_x >= 285 & pix_x <=300 & pix_y >= 253 & pix_y <=253 ) | (pix_x >= 375 & pix_x <=466 & pix_y >= 253 & pix_y <=253 ) | (pix_x >= 287 & pix_x <=299 & pix_y >= 254 & pix_y <=254 ) | (pix_x >= 376 & pix_x <=466 & pix_y >= 254 & pix_y <=254 ) | (pix_x >= 289 & pix_x <=298 & pix_y >= 255 & pix_y <=255 ) | (pix_x >= 378 & pix_x <=466 & pix_y >= 255 & pix_y <=255 ) | (pix_x >= 382 & pix_x <=466 & pix_y >= 256 & pix_y <=256 ) | (pix_x >= 383 & pix_x <=466 & pix_y >= 257 & pix_y <=257 ) | (pix_x >= 383 & pix_x <=466 & pix_y >= 258 & pix_y <=258 ) | (pix_x >= 384 & pix_x <=466 & pix_y >= 259 & pix_y <=258 ) | (pix_x >= 386 & pix_x <=434 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 437 & pix_x <=466 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 386 & pix_x <=430 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 438 & pix_x <=466 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 387 & pix_x <=428 & pix_y >= 261 & pix_y <=261 ) | (pix_x >= 439 & pix_x <=466 & pix_y >= 261 & pix_y <=261 ) | (pix_x >= 388 & pix_x <=427 & pix_y >= 262 & pix_y <=262 ) | (pix_x >= 439 & pix_x <=466 & pix_y >= 262 & pix_y <=262 ) | (pix_x >= 390 & pix_x <=427 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 439 & pix_x <=466 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 385 & pix_x <=424 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 437 & pix_x <=467 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 385 & pix_x <=420 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 437 & pix_x <=440 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 445 & pix_x <=467 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 385 & pix_x <=420 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 445 & pix_x <=466 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 392 & pix_x <=419 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 445 & pix_x <=465 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 393 & pix_x <=420 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 445 & pix_x <=465 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 394 & pix_x <=420 & pix_y >= 269 & pix_y <=269 ) | (pix_x >= 446 & pix_x <=464 & pix_y >= 269 & pix_y <=269 ) | (pix_x >= 394 & pix_x <=420 & pix_y >= 270 & pix_y <=270 ) | (pix_x >= 446 & pix_x <=464 & pix_y >= 270 & pix_y <=270 ) | (pix_x >= 394 & pix_x <=421 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 433 & pix_x <=464 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 393 & pix_x <=424 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 429 & pix_x <=463 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 393 & pix_x <=456 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 460 & pix_x <=462 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 394 & pix_x <=455 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 395 & pix_x <=459 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 395 & pix_x <=460 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 396 & pix_x <=460 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 396 & pix_x <=460 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 396 & pix_x <=460 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 396 & pix_x <=460 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 396 & pix_x <=459 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 396 & pix_x <=459 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 396 & pix_x <=432 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 441 & pix_x <=458 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 396 & pix_x <=435 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 441 & pix_x <=458 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 396 & pix_x <=440 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 444 & pix_x <=457 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 396 & pix_x <=440 & pix_y >= 286 & pix_y <=286 ) | (pix_x >= 448 & pix_x <=456 & pix_y >= 286 & pix_y <=286 ) | (pix_x >= 396 & pix_x <=436 & pix_y >= 287 & pix_y <=287 ) | (pix_x >= 454 & pix_x <=456 & pix_y >= 287 & pix_y <=287 ) | (pix_x >= 396 & pix_x <=429 & pix_y >= 288 & pix_y <=288 ) | (pix_x >= 396 & pix_x <=430 & pix_y >= 289 & pix_y <=289 ) | (pix_x >= 397 & pix_x <=432 & pix_y >= 290 & pix_y <=290 ) | (pix_x >= 397 & pix_x <=436 & pix_y >= 291 & pix_y <=291 ) | (pix_x >= 397 & pix_x <=443 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 449 & pix_x <=443 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 398 & pix_x <=445 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 448 & pix_x <=449 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 398 & pix_x <=449 & pix_y >= 294 & pix_y <=294 ) | (pix_x >= 398 & pix_x <=448 & pix_y >= 295 & pix_y <=295 ) | (pix_x >= 401 & pix_x <=448 & pix_y >= 296 & pix_y <=296 ) | (pix_x >= 401 & pix_x <=448 & pix_y >= 297 & pix_y <=297 ) | (pix_x >= 401 & pix_x <=448 & pix_y >= 298 & pix_y <=298 ) | (pix_x >= 403 & pix_x <=448 & pix_y >= 299 & pix_y <=299 ) | (pix_x >= 405 & pix_x <=448 & pix_y >= 300 & pix_y <=300 ) | (pix_x >= 406 & pix_x <=448 & pix_y >= 301 & pix_y <=301 ) | (pix_x >= 408 & pix_x <=448 & pix_y >= 302 & pix_y <=302 ) | (pix_x >= 409 & pix_x <=448 & pix_y >= 303 & pix_y <=303 ) | (pix_x >= 412 & pix_x <=448 & pix_y >= 304 & pix_y <=304 ) | (pix_x >= 412 & pix_x <=448 & pix_y >= 305 & pix_y <=305 ) | (pix_x >= 413 & pix_x <=448 & pix_y >= 306 & pix_y <=306 ) | (pix_x >= 415 & pix_x <=448 & pix_y >= 307 & pix_y <=307 ) | (pix_x >= 418 & pix_x <=448 & pix_y >= 308 & pix_y <=308 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 309 & pix_y <=309 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 310 & pix_y <=310 ) | (pix_x >= 421 & pix_x <=448 & pix_y >= 311 & pix_y <=311 ) | (pix_x >= 421 & pix_x <=448 & pix_y >= 312 & pix_y <=312 ) | (pix_x >= 423 & pix_x <=447 & pix_y >= 313 & pix_y <=313 ) | (pix_x >= 425 & pix_x <=447 & pix_y >= 314 & pix_y <=314 ) | (pix_x >= 428 & pix_x <=446 & pix_y >= 315 & pix_y <=315 ) | (pix_x >= 430 & pix_x <=446 & pix_y >= 316 & pix_y <=316 ) | (pix_x >= 435 & pix_x <=445 & pix_y >= 317 & pix_y <=317 ) | (pix_x >= 436 & pix_x <=444 & pix_y >= 318 & pix_y <=318 ) | (pix_x >= 437 & pix_x <=444 & pix_y >= 319 & pix_y <=319 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 320 & pix_y <=319 ) | (pix_x >= 288 & pix_x <=444 & pix_y >= 348 & pix_y <=319 ) | (pix_x >= 297 & pix_x <=305 & pix_y >= 348 & pix_y <=348 ) | (pix_x >= 287 & pix_x <=288 & pix_y >= 349 & pix_y <=349 ) | (pix_x >= 297 & pix_x <=307 & pix_y >= 349 & pix_y <=349 ) | (pix_x >= 287 & pix_x <=288 & pix_y >= 350 & pix_y <=350 ) | (pix_x >= 297 & pix_x <=308 & pix_y >= 350 & pix_y <=350 ) | (pix_x >= 286 & pix_x <=288 & pix_y >= 351 & pix_y <=351 ) | (pix_x >= 297 & pix_x <=308 & pix_y >= 351 & pix_y <=351 ) | (pix_x >= 290 & pix_x <=312 & pix_y >= 352 & pix_y <=352 ) | (pix_x >= 289 & pix_x <=312 & pix_y >= 353 & pix_y <=353 ) | (pix_x >= 289 & pix_x <=312 & pix_y >= 354 & pix_y <=354 ) | (pix_x >= 289 & pix_x <=314 & pix_y >= 355 & pix_y <=355 ) | (pix_x >= 289 & pix_x <=315 & pix_y >= 356 & pix_y <=356 ) | (pix_x >= 353 & pix_x <=315 & pix_y >= 356 & pix_y <=356 ) | (pix_x >= 289 & pix_x <=314 & pix_y >= 357 & pix_y <=357 ) | (pix_x >= 353 & pix_x <=314 & pix_y >= 357 & pix_y <=357 ) | (pix_x >= 289 & pix_x <=313 & pix_y >= 358 & pix_y <=358 ) | (pix_x >= 350 & pix_x <=353 & pix_y >= 358 & pix_y <=358 ) | (pix_x >= 289 & pix_x <=312 & pix_y >= 359 & pix_y <=359 ) | (pix_x >= 350 & pix_x <=353 & pix_y >= 359 & pix_y <=359 ) | (pix_x >= 285 & pix_x <=312 & pix_y >= 360 & pix_y <=360 ) | (pix_x >= 326 & pix_x <=328 & pix_y >= 360 & pix_y <=360 ) | (pix_x >= 337 & pix_x <=338 & pix_y >= 360 & pix_y <=360 ) | (pix_x >= 346 & pix_x <=352 & pix_y >= 360 & pix_y <=360 ) | (pix_x >= 285 & pix_x <=312 & pix_y >= 361 & pix_y <=361 ) | (pix_x >= 324 & pix_x <=336 & pix_y >= 361 & pix_y <=361 ) | (pix_x >= 345 & pix_x <=352 & pix_y >= 361 & pix_y <=361 ) | (pix_x >= 285 & pix_x <=312 & pix_y >= 362 & pix_y <=362 ) | (pix_x >= 323 & pix_x <=336 & pix_y >= 362 & pix_y <=362 ) | (pix_x >= 343 & pix_x <=352 & pix_y >= 362 & pix_y <=362 ) | (pix_x >= 285 & pix_x <=312 & pix_y >= 363 & pix_y <=363 ) | (pix_x >= 322 & pix_x <=336 & pix_y >= 363 & pix_y <=363 ) | (pix_x >= 340 & pix_x <=351 & pix_y >= 363 & pix_y <=363 ) | (pix_x >= 285 & pix_x <=311 & pix_y >= 364 & pix_y <=364 ) | (pix_x >= 321 & pix_x <=350 & pix_y >= 364 & pix_y <=364 ) | (pix_x >= 285 & pix_x <=310 & pix_y >= 365 & pix_y <=365 ) | (pix_x >= 321 & pix_x <=350 & pix_y >= 365 & pix_y <=365 ) | (pix_x >= 285 & pix_x <=310 & pix_y >= 366 & pix_y <=366 ) | (pix_x >= 321 & pix_x <=350 & pix_y >= 366 & pix_y <=366 ) | (pix_x >= 285 & pix_x <=309 & pix_y >= 367 & pix_y <=367 ) | (pix_x >= 321 & pix_x <=349 & pix_y >= 367 & pix_y <=367 ) | (pix_x >= 285 & pix_x <=308 & pix_y >= 368 & pix_y <=368 ) | (pix_x >= 317 & pix_x <=349 & pix_y >= 368 & pix_y <=368 ) | (pix_x >= 285 & pix_x <=308 & pix_y >= 369 & pix_y <=369 ) | (pix_x >= 317 & pix_x <=348 & pix_y >= 369 & pix_y <=369 ) | (pix_x >= 286 & pix_x <=307 & pix_y >= 370 & pix_y <=370 ) | (pix_x >= 317 & pix_x <=347 & pix_y >= 370 & pix_y <=370 ) | (pix_x >= 288 & pix_x <=304 & pix_y >= 371 & pix_y <=371 ) | (pix_x >= 317 & pix_x <=347 & pix_y >= 371 & pix_y <=371 ) | (pix_x >= 291 & pix_x <=302 & pix_y >= 372 & pix_y <=372 ) | (pix_x >= 317 & pix_x <=346 & pix_y >= 372 & pix_y <=372 ) | (pix_x >= 424 & pix_x <=346 & pix_y >= 372 & pix_y <=372 ) | (pix_x >= 292 & pix_x <=299 & pix_y >= 373 & pix_y <=373 ) | (pix_x >= 317 & pix_x <=345 & pix_y >= 373 & pix_y <=373 ) | (pix_x >= 424 & pix_x <=345 & pix_y >= 373 & pix_y <=373 ) | (pix_x >= 268 & pix_x <=345 & pix_y >= 374 & pix_y <=373 ) | (pix_x >= 293 & pix_x <=297 & pix_y >= 374 & pix_y <=374 ) | (pix_x >= 317 & pix_x <=344 & pix_y >= 374 & pix_y <=374 ) | (pix_x >= 425 & pix_x <=344 & pix_y >= 374 & pix_y <=374 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 375 & pix_y <=375 ) | (pix_x >= 293 & pix_x <=296 & pix_y >= 375 & pix_y <=375 ) | (pix_x >= 317 & pix_x <=344 & pix_y >= 375 & pix_y <=375 ) | (pix_x >= 425 & pix_x <=344 & pix_y >= 375 & pix_y <=375 ) | (pix_x >= 268 & pix_x <=344 & pix_y >= 376 & pix_y <=375 ) | (pix_x >= 272 & pix_x <=344 & pix_y >= 376 & pix_y <=375 ) | (pix_x >= 293 & pix_x <=296 & pix_y >= 376 & pix_y <=376 ) | (pix_x >= 313 & pix_x <=343 & pix_y >= 376 & pix_y <=376 ) | (pix_x >= 425 & pix_x <=343 & pix_y >= 376 & pix_y <=376 ) | (pix_x >= 272 & pix_x <=343 & pix_y >= 377 & pix_y <=376 ) | (pix_x >= 294 & pix_x <=296 & pix_y >= 377 & pix_y <=377 ) | (pix_x >= 313 & pix_x <=342 & pix_y >= 377 & pix_y <=377 ) | (pix_x >= 425 & pix_x <=342 & pix_y >= 377 & pix_y <=377 ) | (pix_x >= 269 & pix_x <=272 & pix_y >= 378 & pix_y <=378 ) | (pix_x >= 313 & pix_x <=341 & pix_y >= 378 & pix_y <=378 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 378 & pix_y <=378 ) | (pix_x >= 269 & pix_x <=272 & pix_y >= 379 & pix_y <=379 ) | (pix_x >= 313 & pix_x <=340 & pix_y >= 379 & pix_y <=379 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 379 & pix_y <=379 ) | (pix_x >= 269 & pix_x <=272 & pix_y >= 380 & pix_y <=380 ) | (pix_x >= 313 & pix_x <=340 & pix_y >= 380 & pix_y <=380 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 380 & pix_y <=380 ) | (pix_x >= 269 & pix_x <=273 & pix_y >= 381 & pix_y <=381 ) | (pix_x >= 289 & pix_x <=273 & pix_y >= 381 & pix_y <=381 ) | (pix_x >= 313 & pix_x <=339 & pix_y >= 381 & pix_y <=381 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 381 & pix_y <=381 ) | (pix_x >= 269 & pix_x <=274 & pix_y >= 382 & pix_y <=382 ) | (pix_x >= 289 & pix_x <=274 & pix_y >= 382 & pix_y <=382 ) | (pix_x >= 313 & pix_x <=338 & pix_y >= 382 & pix_y <=382 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 382 & pix_y <=382 ) | (pix_x >= 269 & pix_x <=274 & pix_y >= 383 & pix_y <=383 ) | (pix_x >= 289 & pix_x <=274 & pix_y >= 383 & pix_y <=383 ) | (pix_x >= 313 & pix_x <=337 & pix_y >= 383 & pix_y <=383 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 383 & pix_y <=383 ) | (pix_x >= 269 & pix_x <=280 & pix_y >= 384 & pix_y <=384 ) | (pix_x >= 285 & pix_x <=288 & pix_y >= 384 & pix_y <=384 ) | (pix_x >= 317 & pix_x <=336 & pix_y >= 384 & pix_y <=384 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 384 & pix_y <=384 ) | (pix_x >= 269 & pix_x <=280 & pix_y >= 385 & pix_y <=385 ) | (pix_x >= 317 & pix_x <=336 & pix_y >= 385 & pix_y <=385 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 385 & pix_y <=385 ) | (pix_x >= 270 & pix_x <=279 & pix_y >= 386 & pix_y <=386 ) | (pix_x >= 316 & pix_x <=336 & pix_y >= 386 & pix_y <=386 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 386 & pix_y <=386 ) | (pix_x >= 270 & pix_x <=279 & pix_y >= 387 & pix_y <=387 ) | (pix_x >= 315 & pix_x <=336 & pix_y >= 387 & pix_y <=387 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 387 & pix_y <=387 ) | (pix_x >= 270 & pix_x <=282 & pix_y >= 388 & pix_y <=388 ) | (pix_x >= 305 & pix_x <=336 & pix_y >= 388 & pix_y <=388 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 388 & pix_y <=388 ) | (pix_x >= 271 & pix_x <=284 & pix_y >= 389 & pix_y <=389 ) | (pix_x >= 304 & pix_x <=335 & pix_y >= 389 & pix_y <=389 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 389 & pix_y <=389 ) | (pix_x >= 271 & pix_x <=286 & pix_y >= 390 & pix_y <=390 ) | (pix_x >= 302 & pix_x <=334 & pix_y >= 390 & pix_y <=390 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 390 & pix_y <=390 ) | (pix_x >= 271 & pix_x <=287 & pix_y >= 391 & pix_y <=391 ) | (pix_x >= 301 & pix_x <=334 & pix_y >= 391 & pix_y <=391 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 391 & pix_y <=391 ) | (pix_x >= 272 & pix_x <=290 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 300 & pix_x <=333 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 272 & pix_x <=294 & pix_y >= 393 & pix_y <=393 ) | (pix_x >= 297 & pix_x <=333 & pix_y >= 393 & pix_y <=393 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 393 & pix_y <=393 ) | (pix_x >= 272 & pix_x <=333 & pix_y >= 394 & pix_y <=394 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 394 & pix_y <=394 ) | (pix_x >= 273 & pix_x <=332 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 273 & pix_x <=332 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 273 & pix_x <=331 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 273 & pix_x <=331 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 274 & pix_x <=331 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 275 & pix_x <=331 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 276 & pix_x <=330 & pix_y >= 403 & pix_y <=403 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 403 & pix_y <=403 ) | (pix_x >= 276 & pix_x <=329 & pix_y >= 404 & pix_y <=404 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 404 & pix_y <=404 ) | (pix_x >= 276 & pix_x <=329 & pix_y >= 405 & pix_y <=405 ) | (pix_x >= 427 & pix_x <=430 & pix_y >= 405 & pix_y <=405 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 406 & pix_y <=406 ) | (pix_x >= 427 & pix_x <=430 & pix_y >= 406 & pix_y <=406 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 407 & pix_y <=407 ) | (pix_x >= 427 & pix_x <=430 & pix_y >= 407 & pix_y <=407 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 408 & pix_y <=408 ) | (pix_x >= 427 & pix_x <=428 & pix_y >= 408 & pix_y <=408 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 409 & pix_y <=409 ) | (pix_x >= 427 & pix_x <=428 & pix_y >= 409 & pix_y <=409 ) | (pix_x >= 279 & pix_x <=328 & pix_y >= 410 & pix_y <=410 ) | (pix_x >= 426 & pix_x <=427 & pix_y >= 410 & pix_y <=410 ) | (pix_x >= 429 & pix_x <=430 & pix_y >= 410 & pix_y <=410 ) | (pix_x >= 279 & pix_x <=328 & pix_y >= 411 & pix_y <=411 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 411 & pix_y <=411 ) | (pix_x >= 279 & pix_x <=328 & pix_y >= 412 & pix_y <=412 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 412 & pix_y <=412 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 413 & pix_y <=413 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 413 & pix_y <=413 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 281 & pix_x <=327 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 281 & pix_x <=327 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 281 & pix_x <=327 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 283 & pix_x <=326 & pix_y >= 420 & pix_y <=420 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 420 & pix_y <=420 ) | (pix_x >= 283 & pix_x <=325 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 425 & pix_x <=431 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 424 & pix_y <=424 ) | (pix_x >= 426 & pix_x <=430 & pix_y >= 424 & pix_y <=424 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 425 & pix_y <=425 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 425 & pix_y <=425 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 286 & pix_x <=323 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 286 & pix_x <=323 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 425 & pix_x <=431 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 287 & pix_x <=322 & pix_y >= 429 & pix_y <=429 ) | (pix_x >= 424 & pix_x <=425 & pix_y >= 429 & pix_y <=429 ) | (pix_x >= 427 & pix_x <=430 & pix_y >= 429 & pix_y <=429 ) | (pix_x >= 287 & pix_x <=322 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 423 & pix_x <=426 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 429 & pix_x <=430 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 288 & pix_x <=321 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 423 & pix_x <=430 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 289 & pix_x <=320 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 423 & pix_x <=430 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 289 & pix_x <=320 & pix_y >= 433 & pix_y <=433 ) | (pix_x >= 423 & pix_x <=430 & pix_y >= 433 & pix_y <=433 ) | (pix_x >= 289 & pix_x <=320 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 423 & pix_x <=425 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 429 & pix_x <=431 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 290 & pix_x <=319 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 422 & pix_x <=430 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 291 & pix_x <=318 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 422 & pix_x <=430 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 291 & pix_x <=317 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 424 & pix_x <=430 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 291 & pix_x <=316 & pix_y >= 438 & pix_y <=438 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 438 & pix_y <=438 ) | (pix_x >= 429 & pix_x <=430 & pix_y >= 438 & pix_y <=438 ) | (pix_x >= 292 & pix_x <=316 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 421 & pix_x <=424 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 428 & pix_x <=429 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 432 & pix_x <=429 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 292 & pix_x <=315 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 420 & pix_x <=427 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 430 & pix_x <=432 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 293 & pix_x <=314 & pix_y >= 441 & pix_y <=441 ) | (pix_x >= 421 & pix_x <=428 & pix_y >= 441 & pix_y <=441 ) | (pix_x >= 294 & pix_x <=314 & pix_y >= 442 & pix_y <=442 ) | (pix_x >= 421 & pix_x <=423 & pix_y >= 442 & pix_y <=442 ) | (pix_x >= 425 & pix_x <=430 & pix_y >= 442 & pix_y <=442 ) | (pix_x >= 294 & pix_x <=313 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 419 & pix_x <=313 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 421 & pix_x <=423 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 428 & pix_x <=431 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 294 & pix_x <=313 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 419 & pix_x <=313 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 421 & pix_x <=425 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 429 & pix_x <=432 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 295 & pix_x <=312 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 422 & pix_x <=427 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 295 & pix_x <=311 & pix_y >= 446 & pix_y <=446 ) | (pix_x >= 421 & pix_x <=430 & pix_y >= 446 & pix_y <=446 ) | (pix_x >= 296 & pix_x <=311 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 420 & pix_x <=422 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 428 & pix_x <=431 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 297 & pix_x <=310 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 420 & pix_x <=423 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 297 & pix_x <=309 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 417 & pix_x <=309 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 421 & pix_x <=424 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 298 & pix_x <=309 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 421 & pix_x <=424 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 299 & pix_x <=308 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 419 & pix_x <=422 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 299 & pix_x <=308 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 419 & pix_x <=422 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 300 & pix_x <=307 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 420 & pix_x <=424 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 300 & pix_x <=306 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 420 & pix_x <=424 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 301 & pix_x <=306 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 419 & pix_x <=421 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 303 & pix_x <=304 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=427 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 433 & pix_x <=427 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 304 & pix_x <=427 & pix_y >= 457 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=427 & pix_y >= 457 & pix_y <=457 ) | (pix_x >= 433 & pix_x <=427 & pix_y >= 457 & pix_y <=457 ) | (pix_x >= 419 & pix_x <=427 & pix_y >= 458 & pix_y <=458 ) | (pix_x >= 433 & pix_x <=427 & pix_y >= 458 & pix_y <=458 ) | (pix_x >= 420 & pix_x <=421 & pix_y >= 459 & pix_y <=459 ) | (pix_x >= 426 & pix_x <=427 & pix_y >= 459 & pix_y <=459 ) | (pix_x >= 433 & pix_x <=427 & pix_y >= 459 & pix_y <=459 ) | (pix_x >= 418 & pix_x <=420 & pix_y >= 460 & pix_y <=460 ) | (pix_x >= 433 & pix_x <=420 & pix_y >= 460 & pix_y <=460 ) | (pix_x >= 417 & pix_x <=420 & pix_y >= 461 & pix_y <=461 ) | (pix_x >= 433 & pix_x <=420 & pix_y >= 461 & pix_y <=461 ) | (pix_x >= 417 & pix_x <=421 & pix_y >= 462 & pix_y <=462 ) | (pix_x >= 433 & pix_x <=421 & pix_y >= 462 & pix_y <=462 ) | (pix_x >= 419 & pix_x <=421 & pix_y >= 463 & pix_y <=463 ) | (pix_x >= 433 & pix_x <=421 & pix_y >= 463 & pix_y <=463 ) | (pix_x >= 413 & pix_x <=421 & pix_y >= 464 & pix_y <=463 ) | (pix_x >= 417 & pix_x <=419 & pix_y >= 464 & pix_y <=464 ) | (pix_x >= 413 & pix_x <=419 & pix_y >= 465 & pix_y <=464 ) | (pix_x >= 417 & pix_x <=419 & pix_y >= 465 & pix_y <=465 ) | (pix_x >= 417 & pix_x <=420 & pix_y >= 466 & pix_y <=466 ) | (pix_x >= 417 & pix_x <=420 & pix_y >= 467 & pix_y <=467 ) | (pix_x >= 417 & pix_x <=419 & pix_y >= 468 & pix_y <=468 ) | (pix_x >= 416 & pix_x <=418 & pix_y >= 470 & pix_y <=470 ) | (pix_x >= 424 & pix_x <=418 & pix_y >= 470 & pix_y <=470 ) | (pix_x >= 416 & pix_x <=419 & pix_y >= 471 & pix_y <=471 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 471 & pix_y <=471 ) | (pix_x >= 417 & pix_x <=424 & pix_y >= 472 & pix_y <=472 ) ;


//---------GREEN---------


assign g_out =  (pix_x >= 406 & pix_x <=411 & pix_y >= 113 & pix_y <=113 ) | (pix_x >= 417 & pix_x <=420 & pix_y >= 113 & pix_y <=113 ) | (pix_x >= 393 & pix_x <=425 & pix_y >= 114 & pix_y <=114 ) | (pix_x >= 390 & pix_x <=427 & pix_y >= 115 & pix_y <=115 ) | (pix_x >= 389 & pix_x <=427 & pix_y >= 116 & pix_y <=116 ) | (pix_x >= 385 & pix_x <=428 & pix_y >= 117 & pix_y <=117 ) | (pix_x >= 382 & pix_x <=429 & pix_y >= 118 & pix_y <=118 ) | (pix_x >= 381 & pix_x <=430 & pix_y >= 119 & pix_y <=119 ) | (pix_x >= 380 & pix_x <=430 & pix_y >= 120 & pix_y <=120 ) | (pix_x >= 380 & pix_x <=430 & pix_y >= 121 & pix_y <=121 ) | (pix_x >= 378 & pix_x <=432 & pix_y >= 122 & pix_y <=122 ) | (pix_x >= 377 & pix_x <=432 & pix_y >= 123 & pix_y <=123 ) | (pix_x >= 377 & pix_x <=435 & pix_y >= 124 & pix_y <=124 ) | (pix_x >= 378 & pix_x <=435 & pix_y >= 125 & pix_y <=125 ) | (pix_x >= 380 & pix_x <=436 & pix_y >= 126 & pix_y <=126 ) | (pix_x >= 380 & pix_x <=436 & pix_y >= 127 & pix_y <=127 ) | (pix_x >= 381 & pix_x <=436 & pix_y >= 128 & pix_y <=128 ) | (pix_x >= 381 & pix_x <=437 & pix_y >= 129 & pix_y <=129 ) | (pix_x >= 381 & pix_x <=438 & pix_y >= 130 & pix_y <=130 ) | (pix_x >= 381 & pix_x <=440 & pix_y >= 131 & pix_y <=131 ) | (pix_x >= 381 & pix_x <=441 & pix_y >= 132 & pix_y <=132 ) | (pix_x >= 381 & pix_x <=442 & pix_y >= 133 & pix_y <=133 ) | (pix_x >= 381 & pix_x <=444 & pix_y >= 134 & pix_y <=134 ) | (pix_x >= 381 & pix_x <=445 & pix_y >= 135 & pix_y <=135 ) | (pix_x >= 381 & pix_x <=446 & pix_y >= 136 & pix_y <=136 ) | (pix_x >= 381 & pix_x <=447 & pix_y >= 137 & pix_y <=137 ) | (pix_x >= 381 & pix_x <=448 & pix_y >= 138 & pix_y <=138 ) | (pix_x >= 380 & pix_x <=448 & pix_y >= 139 & pix_y <=139 ) | (pix_x >= 380 & pix_x <=449 & pix_y >= 140 & pix_y <=140 ) | (pix_x >= 379 & pix_x <=449 & pix_y >= 141 & pix_y <=141 ) | (pix_x >= 379 & pix_x <=449 & pix_y >= 142 & pix_y <=142 ) | (pix_x >= 379 & pix_x <=450 & pix_y >= 143 & pix_y <=143 ) | (pix_x >= 381 & pix_x <=450 & pix_y >= 144 & pix_y <=144 ) | (pix_x >= 381 & pix_x <=451 & pix_y >= 145 & pix_y <=145 ) | (pix_x >= 380 & pix_x <=451 & pix_y >= 146 & pix_y <=146 ) | (pix_x >= 376 & pix_x <=451 & pix_y >= 147 & pix_y <=146 ) | (pix_x >= 379 & pix_x <=452 & pix_y >= 147 & pix_y <=147 ) | (pix_x >= 374 & pix_x <=452 & pix_y >= 148 & pix_y <=148 ) | (pix_x >= 372 & pix_x <=453 & pix_y >= 149 & pix_y <=149 ) | (pix_x >= 372 & pix_x <=375 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 377 & pix_x <=404 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 407 & pix_x <=454 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 369 & pix_x <=372 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 377 & pix_x <=403 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 409 & pix_x <=454 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 368 & pix_x <=376 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 379 & pix_x <=387 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 390 & pix_x <=402 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 412 & pix_x <=455 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 379 & pix_x <=396 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 410 & pix_x <=455 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 379 & pix_x <=390 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 408 & pix_x <=456 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 380 & pix_x <=381 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 387 & pix_x <=388 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 406 & pix_x <=412 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 416 & pix_x <=456 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 405 & pix_x <=409 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 414 & pix_x <=420 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 422 & pix_x <=457 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 413 & pix_x <=420 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 423 & pix_x <=457 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 409 & pix_x <=416 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 418 & pix_x <=419 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 424 & pix_x <=419 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 427 & pix_x <=457 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 409 & pix_x <=415 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 433 & pix_x <=458 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 360 & pix_x <=458 & pix_y >= 160 & pix_y <=159 ) | (pix_x >= 406 & pix_x <=418 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 433 & pix_x <=458 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 405 & pix_x <=419 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 439 & pix_x <=458 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 405 & pix_x <=418 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 403 & pix_x <=418 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 401 & pix_x <=420 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 401 & pix_x <=421 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 405 & pix_x <=422 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 409 & pix_x <=429 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 410 & pix_x <=435 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 410 & pix_x <=426 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 428 & pix_x <=431 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 433 & pix_x <=440 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 446 & pix_x <=459 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 410 & pix_x <=431 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 436 & pix_x <=441 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 446 & pix_x <=459 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 441 & pix_x <=443 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 446 & pix_x <=459 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 353 & pix_x <=356 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 445 & pix_x <=458 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 410 & pix_x <=417 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 420 & pix_x <=432 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 447 & pix_x <=456 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 411 & pix_x <=416 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 448 & pix_x <=456 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 412 & pix_x <=432 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 449 & pix_x <=456 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 414 & pix_x <=424 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 444 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 450 & pix_x <=455 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 414 & pix_x <=432 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 451 & pix_x <=455 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 422 & pix_x <=432 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 453 & pix_x <=455 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 454 & pix_x <=446 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 423 & pix_x <=431 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 359 & pix_x <=377 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 415 & pix_x <=416 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 423 & pix_x <=431 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 353 & pix_x <=378 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 422 & pix_x <=432 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 457 & pix_x <=448 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 350 & pix_x <=381 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 456 & pix_x <=458 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 352 & pix_x <=384 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 352 & pix_x <=384 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 407 & pix_x <=408 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 457 & pix_x <=459 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 465 & pix_x <=467 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 352 & pix_x <=383 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 424 & pix_x <=417 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 457 & pix_x <=459 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 463 & pix_x <=468 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 352 & pix_x <=384 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 404 & pix_x <=408 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 424 & pix_x <=417 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 457 & pix_x <=458 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 463 & pix_x <=464 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 353 & pix_x <=384 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 403 & pix_x <=408 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 424 & pix_x <=417 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 463 & pix_x <=465 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 356 & pix_x <=384 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 358 & pix_x <=387 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 416 & pix_x <=418 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 462 & pix_x <=465 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 360 & pix_x <=388 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 416 & pix_x <=417 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 454 & pix_x <=455 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 361 & pix_x <=392 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 403 & pix_x <=408 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 442 & pix_x <=445 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 454 & pix_x <=456 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 361 & pix_x <=392 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 403 & pix_x <=408 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 415 & pix_x <=419 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 421 & pix_x <=422 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 442 & pix_x <=445 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 454 & pix_x <=457 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 363 & pix_x <=392 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 403 & pix_x <=408 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 416 & pix_x <=422 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 425 & pix_x <=433 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 442 & pix_x <=444 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 454 & pix_x <=458 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 364 & pix_x <=395 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 403 & pix_x <=408 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 416 & pix_x <=422 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 425 & pix_x <=434 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 442 & pix_x <=444 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 454 & pix_x <=460 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 365 & pix_x <=408 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 416 & pix_x <=437 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 454 & pix_x <=466 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 366 & pix_x <=408 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 416 & pix_x <=437 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 367 & pix_x <=408 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 416 & pix_x <=437 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 445 & pix_x <=446 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 368 & pix_x <=409 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 416 & pix_x <=437 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 445 & pix_x <=446 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 448 & pix_x <=446 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 369 & pix_x <=409 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 441 & pix_x <=446 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 370 & pix_x <=409 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 444 & pix_x <=446 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 453 & pix_x <=467 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 371 & pix_x <=409 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 445 & pix_x <=442 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 453 & pix_x <=454 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 456 & pix_x <=468 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 372 & pix_x <=409 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 441 & pix_x <=443 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 452 & pix_x <=454 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 456 & pix_x <=469 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 373 & pix_x <=409 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 452 & pix_x <=454 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 457 & pix_x <=470 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 374 & pix_x <=409 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 452 & pix_x <=454 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 457 & pix_x <=471 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 374 & pix_x <=409 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 452 & pix_x <=455 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 457 & pix_x <=472 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 375 & pix_x <=409 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 451 & pix_x <=472 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 377 & pix_x <=409 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 452 & pix_x <=474 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 378 & pix_x <=409 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 451 & pix_x <=474 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 378 & pix_x <=409 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 451 & pix_x <=475 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 257 & pix_x <=258 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 268 & pix_x <=258 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 379 & pix_x <=410 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 451 & pix_x <=454 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 456 & pix_x <=476 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 258 & pix_x <=476 & pix_y >= 212 & pix_y <=211 ) | (pix_x >= 268 & pix_x <=476 & pix_y >= 212 & pix_y <=211 ) | (pix_x >= 380 & pix_x <=410 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 450 & pix_x <=453 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 456 & pix_x <=477 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 258 & pix_x <=477 & pix_y >= 213 & pix_y <=212 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 381 & pix_x <=411 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 418 & pix_x <=439 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 450 & pix_x <=478 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 258 & pix_x <=259 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 381 & pix_x <=411 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 419 & pix_x <=439 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 450 & pix_x <=479 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 258 & pix_x <=259 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 382 & pix_x <=411 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 420 & pix_x <=439 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 450 & pix_x <=463 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 465 & pix_x <=480 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 259 & pix_x <=480 & pix_y >= 216 & pix_y <=215 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 383 & pix_x <=413 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 421 & pix_x <=439 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 449 & pix_x <=461 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 465 & pix_x <=481 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 259 & pix_x <=481 & pix_y >= 217 & pix_y <=216 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 383 & pix_x <=414 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 422 & pix_x <=439 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 448 & pix_x <=462 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 465 & pix_x <=481 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 259 & pix_x <=260 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 384 & pix_x <=416 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 424 & pix_x <=438 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 449 & pix_x <=482 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 259 & pix_x <=260 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 269 & pix_x <=271 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 384 & pix_x <=418 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 427 & pix_x <=438 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 449 & pix_x <=483 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 260 & pix_x <=483 & pix_y >= 220 & pix_y <=219 ) | (pix_x >= 270 & pix_x <=271 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 385 & pix_x <=419 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 428 & pix_x <=439 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 441 & pix_x <=439 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 449 & pix_x <=483 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 261 & pix_x <=483 & pix_y >= 221 & pix_y <=220 ) | (pix_x >= 270 & pix_x <=272 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 386 & pix_x <=421 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 432 & pix_x <=440 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 448 & pix_x <=484 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 261 & pix_x <=484 & pix_y >= 222 & pix_y <=221 ) | (pix_x >= 271 & pix_x <=272 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 387 & pix_x <=424 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 448 & pix_x <=484 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 261 & pix_x <=262 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 272 & pix_x <=273 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 387 & pix_x <=429 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 449 & pix_x <=485 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 262 & pix_x <=485 & pix_y >= 224 & pix_y <=223 ) | (pix_x >= 273 & pix_x <=275 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 385 & pix_x <=431 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 451 & pix_x <=485 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 273 & pix_x <=275 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 385 & pix_x <=429 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 452 & pix_x <=485 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 264 & pix_x <=485 & pix_y >= 226 & pix_y <=225 ) | (pix_x >= 274 & pix_x <=276 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 385 & pix_x <=427 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 454 & pix_x <=485 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 264 & pix_x <=485 & pix_y >= 227 & pix_y <=226 ) | (pix_x >= 275 & pix_x <=277 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 385 & pix_x <=426 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 264 & pix_x <=265 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 276 & pix_x <=277 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 385 & pix_x <=424 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 265 & pix_x <=266 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 385 & pix_x <=425 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 429 & pix_x <=435 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 265 & pix_x <=266 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 385 & pix_x <=435 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 456 & pix_x <=470 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 476 & pix_x <=485 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 265 & pix_x <=268 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 385 & pix_x <=435 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 456 & pix_x <=470 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 476 & pix_x <=485 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 266 & pix_x <=270 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 288 & pix_x <=289 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 385 & pix_x <=435 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 455 & pix_x <=465 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 476 & pix_x <=485 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 267 & pix_x <=271 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 288 & pix_x <=290 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 385 & pix_x <=435 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 456 & pix_x <=435 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 458 & pix_x <=461 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 476 & pix_x <=484 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 268 & pix_x <=272 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 289 & pix_x <=293 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 477 & pix_x <=484 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 268 & pix_x <=272 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 290 & pix_x <=293 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 477 & pix_x <=484 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 269 & pix_x <=273 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 292 & pix_x <=293 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 478 & pix_x <=483 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 270 & pix_x <=274 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 481 & pix_x <=483 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 271 & pix_x <=275 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 279 & pix_x <=281 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 481 & pix_x <=482 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 271 & pix_x <=274 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 278 & pix_x <=282 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 385 & pix_x <=436 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 481 & pix_x <=482 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 273 & pix_x <=282 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 385 & pix_x <=437 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 454 & pix_x <=456 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 273 & pix_x <=282 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 385 & pix_x <=392 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 394 & pix_x <=437 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 453 & pix_x <=460 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 275 & pix_x <=283 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 385 & pix_x <=392 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 395 & pix_x <=438 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 454 & pix_x <=461 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 275 & pix_x <=283 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 387 & pix_x <=390 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 395 & pix_x <=439 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 457 & pix_x <=461 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 276 & pix_x <=283 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 387 & pix_x <=390 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 396 & pix_x <=442 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 457 & pix_x <=462 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 277 & pix_x <=284 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 387 & pix_x <=390 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 397 & pix_x <=448 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 453 & pix_x <=463 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 277 & pix_x <=284 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 286 & pix_x <=288 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 388 & pix_x <=389 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 397 & pix_x <=464 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 278 & pix_x <=289 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 297 & pix_x <=289 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 388 & pix_x <=389 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 397 & pix_x <=464 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 279 & pix_x <=288 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 290 & pix_x <=292 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 392 & pix_x <=292 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 397 & pix_x <=464 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 466 & pix_x <=467 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 281 & pix_x <=288 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 290 & pix_x <=293 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 398 & pix_x <=467 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 281 & pix_x <=288 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 290 & pix_x <=293 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 398 & pix_x <=466 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 285 & pix_x <=288 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 291 & pix_x <=294 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 398 & pix_x <=466 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 288 & pix_x <=466 & pix_y >= 252 & pix_y <=251 ) | (pix_x >= 398 & pix_x <=466 & pix_y >= 252 & pix_y <=252 ) | (pix_x >= 399 & pix_x <=465 & pix_y >= 253 & pix_y <=253 ) | (pix_x >= 399 & pix_x <=465 & pix_y >= 254 & pix_y <=254 ) | (pix_x >= 399 & pix_x <=464 & pix_y >= 255 & pix_y <=255 ) | (pix_x >= 399 & pix_x <=465 & pix_y >= 256 & pix_y <=256 ) | (pix_x >= 399 & pix_x <=465 & pix_y >= 257 & pix_y <=257 ) | (pix_x >= 400 & pix_x <=432 & pix_y >= 258 & pix_y <=258 ) | (pix_x >= 438 & pix_x <=465 & pix_y >= 258 & pix_y <=258 ) | (pix_x >= 401 & pix_x <=429 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 439 & pix_x <=465 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 401 & pix_x <=427 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 403 & pix_x <=424 & pix_y >= 261 & pix_y <=261 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 261 & pix_y <=261 ) | (pix_x >= 404 & pix_x <=418 & pix_y >= 262 & pix_y <=262 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 262 & pix_y <=262 ) | (pix_x >= 404 & pix_x <=416 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 440 & pix_x <=453 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 457 & pix_x <=465 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 408 & pix_x <=416 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 441 & pix_x <=416 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 453 & pix_x <=457 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 460 & pix_x <=467 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 408 & pix_x <=414 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 452 & pix_x <=458 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 461 & pix_x <=466 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 408 & pix_x <=411 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 408 & pix_x <=466 & pix_y >= 267 & pix_y <=266 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 463 & pix_x <=465 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 408 & pix_x <=465 & pix_y >= 268 & pix_y <=267 ) | (pix_x >= 449 & pix_x <=465 & pix_y >= 268 & pix_y <=267 ) | (pix_x >= 454 & pix_x <=460 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 463 & pix_x <=465 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 408 & pix_x <=465 & pix_y >= 269 & pix_y <=268 ) | (pix_x >= 456 & pix_x <=465 & pix_y >= 269 & pix_y <=268 ) | (pix_x >= 458 & pix_x <=464 & pix_y >= 269 & pix_y <=269 ) | (pix_x >= 408 & pix_x <=464 & pix_y >= 270 & pix_y <=269 ) | (pix_x >= 457 & pix_x <=464 & pix_y >= 270 & pix_y <=269 ) | (pix_x >= 461 & pix_x <=464 & pix_y >= 270 & pix_y <=270 ) | (pix_x >= 408 & pix_x <=411 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 457 & pix_x <=411 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 462 & pix_x <=464 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 407 & pix_x <=410 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 432 & pix_x <=448 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 461 & pix_x <=462 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 407 & pix_x <=410 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 416 & pix_x <=424 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 433 & pix_x <=434 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 436 & pix_x <=451 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 407 & pix_x <=410 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 415 & pix_x <=429 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 439 & pix_x <=453 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 407 & pix_x <=433 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 441 & pix_x <=456 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 407 & pix_x <=436 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 407 & pix_x <=428 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 430 & pix_x <=437 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 445 & pix_x <=460 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 407 & pix_x <=427 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 433 & pix_x <=440 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 447 & pix_x <=460 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 407 & pix_x <=426 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 435 & pix_x <=440 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 437 & pix_x <=441 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 438 & pix_x <=442 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 451 & pix_x <=459 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 445 & pix_x <=427 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 453 & pix_x <=458 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 445 & pix_x <=457 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 447 & pix_x <=456 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 406 & pix_x <=427 & pix_y >= 286 & pix_y <=286 ) | (pix_x >= 456 & pix_x <=427 & pix_y >= 286 & pix_y <=286 ) | (pix_x >= 406 & pix_x <=415 & pix_y >= 287 & pix_y <=287 ) | (pix_x >= 417 & pix_x <=427 & pix_y >= 287 & pix_y <=287 ) | (pix_x >= 411 & pix_x <=424 & pix_y >= 288 & pix_y <=288 ) | (pix_x >= 412 & pix_x <=422 & pix_y >= 289 & pix_y <=289 ) | (pix_x >= 413 & pix_x <=420 & pix_y >= 290 & pix_y <=290 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 291 & pix_y <=291 ) | (pix_x >= 427 & pix_x <=429 & pix_y >= 291 & pix_y <=291 ) | (pix_x >= 415 & pix_x <=416 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 435 & pix_x <=442 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 421 & pix_x <=444 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 449 & pix_x <=444 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 419 & pix_x <=449 & pix_y >= 294 & pix_y <=294 ) | (pix_x >= 417 & pix_x <=448 & pix_y >= 295 & pix_y <=295 ) | (pix_x >= 417 & pix_x <=448 & pix_y >= 296 & pix_y <=296 ) | (pix_x >= 417 & pix_x <=447 & pix_y >= 297 & pix_y <=297 ) | (pix_x >= 417 & pix_x <=447 & pix_y >= 298 & pix_y <=298 ) | (pix_x >= 417 & pix_x <=447 & pix_y >= 299 & pix_y <=299 ) | (pix_x >= 417 & pix_x <=447 & pix_y >= 300 & pix_y <=300 ) | (pix_x >= 417 & pix_x <=447 & pix_y >= 301 & pix_y <=301 ) | (pix_x >= 417 & pix_x <=448 & pix_y >= 302 & pix_y <=302 ) | (pix_x >= 417 & pix_x <=448 & pix_y >= 303 & pix_y <=303 ) | (pix_x >= 419 & pix_x <=448 & pix_y >= 304 & pix_y <=304 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 305 & pix_y <=305 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 306 & pix_y <=306 ) | (pix_x >= 422 & pix_x <=448 & pix_y >= 307 & pix_y <=307 ) | (pix_x >= 423 & pix_x <=448 & pix_y >= 308 & pix_y <=308 ) | (pix_x >= 425 & pix_x <=448 & pix_y >= 309 & pix_y <=309 ) | (pix_x >= 425 & pix_x <=448 & pix_y >= 310 & pix_y <=310 ) | (pix_x >= 425 & pix_x <=442 & pix_y >= 311 & pix_y <=311 ) | (pix_x >= 444 & pix_x <=448 & pix_y >= 311 & pix_y <=311 ) | (pix_x >= 427 & pix_x <=440 & pix_y >= 312 & pix_y <=312 ) | (pix_x >= 445 & pix_x <=447 & pix_y >= 312 & pix_y <=312 ) | (pix_x >= 428 & pix_x <=439 & pix_y >= 313 & pix_y <=313 ) | (pix_x >= 444 & pix_x <=447 & pix_y >= 313 & pix_y <=313 ) | (pix_x >= 435 & pix_x <=438 & pix_y >= 314 & pix_y <=314 ) | (pix_x >= 444 & pix_x <=446 & pix_y >= 314 & pix_y <=314 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 315 & pix_y <=315 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 316 & pix_y <=316 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 317 & pix_y <=317 ) | (pix_x >= 353 & pix_x <=444 & pix_y >= 359 & pix_y <=317 ) | (pix_x >= 351 & pix_x <=352 & pix_y >= 360 & pix_y <=360 ) | (pix_x >= 351 & pix_x <=352 & pix_y >= 361 & pix_y <=361 ) | (pix_x >= 349 & pix_x <=351 & pix_y >= 362 & pix_y <=362 ) | (pix_x >= 347 & pix_x <=350 & pix_y >= 363 & pix_y <=363 ) | (pix_x >= 345 & pix_x <=350 & pix_y >= 364 & pix_y <=364 ) | (pix_x >= 345 & pix_x <=349 & pix_y >= 365 & pix_y <=365 ) | (pix_x >= 341 & pix_x <=345 & pix_y >= 366 & pix_y <=366 ) | (pix_x >= 348 & pix_x <=349 & pix_y >= 366 & pix_y <=366 ) | (pix_x >= 329 & pix_x <=344 & pix_y >= 367 & pix_y <=367 ) | (pix_x >= 348 & pix_x <=349 & pix_y >= 367 & pix_y <=367 ) | (pix_x >= 333 & pix_x <=348 & pix_y >= 368 & pix_y <=368 ) | (pix_x >= 333 & pix_x <=347 & pix_y >= 369 & pix_y <=369 ) | (pix_x >= 334 & pix_x <=347 & pix_y >= 370 & pix_y <=370 ) | (pix_x >= 336 & pix_x <=346 & pix_y >= 371 & pix_y <=371 ) | (pix_x >= 337 & pix_x <=345 & pix_y >= 372 & pix_y <=372 ) | (pix_x >= 337 & pix_x <=345 & pix_y >= 373 & pix_y <=373 ) | (pix_x >= 337 & pix_x <=344 & pix_y >= 374 & pix_y <=374 ) | (pix_x >= 337 & pix_x <=344 & pix_y >= 375 & pix_y <=375 ) | (pix_x >= 337 & pix_x <=342 & pix_y >= 376 & pix_y <=376 ) | (pix_x >= 337 & pix_x <=342 & pix_y >= 377 & pix_y <=376 ) | (pix_x >= 340 & pix_x <=342 & pix_y >= 377 & pix_y <=377 ) | (pix_x >= 337 & pix_x <=342 & pix_y >= 378 & pix_y <=377 ) | (pix_x >= 338 & pix_x <=339 & pix_y >= 380 & pix_y <=380 ) | (pix_x >= 338 & pix_x <=339 & pix_y >= 381 & pix_y <=381 ) | (pix_x >= 337 & pix_x <=339 & pix_y >= 382 & pix_y <=381 ) | (pix_x >= 337 & pix_x <=339 & pix_y >= 383 & pix_y <=381 ) | (pix_x >= 272 & pix_x <=339 & pix_y >= 388 & pix_y <=381 ) | (pix_x >= 272 & pix_x <=273 & pix_y >= 389 & pix_y <=389 ) | (pix_x >= 333 & pix_x <=273 & pix_y >= 389 & pix_y <=389 ) | (pix_x >= 332 & pix_x <=333 & pix_y >= 390 & pix_y <=390 ) | (pix_x >= 332 & pix_x <=333 & pix_y >= 391 & pix_y <=391 ) | (pix_x >= 272 & pix_x <=279 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 329 & pix_x <=279 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 331 & pix_x <=333 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 272 & pix_x <=279 & pix_y >= 393 & pix_y <=393 ) | (pix_x >= 329 & pix_x <=333 & pix_y >= 393 & pix_y <=393 ) | (pix_x >= 273 & pix_x <=280 & pix_y >= 394 & pix_y <=394 ) | (pix_x >= 327 & pix_x <=332 & pix_y >= 394 & pix_y <=394 ) | (pix_x >= 273 & pix_x <=281 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 295 & pix_x <=296 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 325 & pix_x <=332 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 273 & pix_x <=282 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 292 & pix_x <=300 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 322 & pix_x <=331 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 274 & pix_x <=283 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 289 & pix_x <=304 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 319 & pix_x <=331 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 274 & pix_x <=283 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 288 & pix_x <=331 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 275 & pix_x <=284 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 287 & pix_x <=296 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 299 & pix_x <=331 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 276 & pix_x <=329 & pix_y >= 403 & pix_y <=403 ) | (pix_x >= 276 & pix_x <=329 & pix_y >= 404 & pix_y <=404 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 405 & pix_y <=405 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 406 & pix_y <=406 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 407 & pix_y <=407 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 408 & pix_y <=408 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 409 & pix_y <=409 ) | (pix_x >= 279 & pix_x <=328 & pix_y >= 410 & pix_y <=410 ) | (pix_x >= 279 & pix_x <=327 & pix_y >= 411 & pix_y <=411 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 412 & pix_y <=412 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 413 & pix_y <=413 ) | (pix_x >= 281 & pix_x <=327 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 281 & pix_x <=327 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 281 & pix_x <=326 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 283 & pix_x <=326 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 427 & pix_x <=428 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 283 & pix_x <=325 & pix_y >= 420 & pix_y <=420 ) | (pix_x >= 283 & pix_x <=325 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 426 & pix_x <=325 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 424 & pix_y <=424 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 425 & pix_y <=425 ) | (pix_x >= 286 & pix_x <=323 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 286 & pix_x <=323 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 287 & pix_x <=322 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 287 & pix_x <=322 & pix_y >= 429 & pix_y <=429 ) | (pix_x >= 288 & pix_x <=321 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 425 & pix_x <=321 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 288 & pix_x <=321 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 424 & pix_x <=426 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 289 & pix_x <=320 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 289 & pix_x <=320 & pix_y >= 433 & pix_y <=433 ) | (pix_x >= 290 & pix_x <=319 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 424 & pix_x <=319 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 290 & pix_x <=318 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 423 & pix_x <=425 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 291 & pix_x <=317 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 424 & pix_x <=426 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 291 & pix_x <=317 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 425 & pix_x <=317 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 292 & pix_x <=315 & pix_y >= 438 & pix_y <=438 ) | (pix_x >= 292 & pix_x <=315 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 292 & pix_x <=314 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 424 & pix_x <=425 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 293 & pix_x <=314 & pix_y >= 441 & pix_y <=441 ) | (pix_x >= 294 & pix_x <=313 & pix_y >= 442 & pix_y <=442 ) | (pix_x >= 294 & pix_x <=312 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 422 & pix_x <=423 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 294 & pix_x <=311 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 423 & pix_x <=311 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 295 & pix_x <=310 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 296 & pix_x <=310 & pix_y >= 446 & pix_y <=446 ) | (pix_x >= 296 & pix_x <=310 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 297 & pix_x <=309 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 421 & pix_x <=422 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 297 & pix_x <=309 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 422 & pix_x <=424 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 299 & pix_x <=308 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 299 & pix_x <=307 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 300 & pix_x <=307 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 420 & pix_x <=422 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 300 & pix_x <=306 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 421 & pix_x <=423 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 301 & pix_x <=305 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 301 & pix_x <=305 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 303 & pix_x <=304 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=421 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 304 & pix_x <=421 & pix_y >= 457 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=421 & pix_y >= 457 & pix_y <=457 ) | (pix_x >= 421 & pix_x <=422 & pix_y >= 458 & pix_y <=458 ) | (pix_x >= 419 & pix_x <=422 & pix_y >= 461 & pix_y <=458 ) ;


//---------BLUE---------


assign b_out =  (pix_x >= 397 & pix_x <=413 & pix_y >= 114 & pix_y <=114 ) | (pix_x >= 417 & pix_x <=425 & pix_y >= 114 & pix_y <=114 ) | (pix_x >= 395 & pix_x <=426 & pix_y >= 115 & pix_y <=115 ) | (pix_x >= 393 & pix_x <=427 & pix_y >= 116 & pix_y <=116 ) | (pix_x >= 390 & pix_x <=428 & pix_y >= 117 & pix_y <=117 ) | (pix_x >= 385 & pix_x <=429 & pix_y >= 118 & pix_y <=118 ) | (pix_x >= 384 & pix_x <=430 & pix_y >= 119 & pix_y <=119 ) | (pix_x >= 382 & pix_x <=429 & pix_y >= 120 & pix_y <=120 ) | (pix_x >= 382 & pix_x <=430 & pix_y >= 121 & pix_y <=121 ) | (pix_x >= 380 & pix_x <=431 & pix_y >= 122 & pix_y <=122 ) | (pix_x >= 379 & pix_x <=383 & pix_y >= 123 & pix_y <=123 ) | (pix_x >= 385 & pix_x <=432 & pix_y >= 123 & pix_y <=123 ) | (pix_x >= 379 & pix_x <=383 & pix_y >= 124 & pix_y <=124 ) | (pix_x >= 385 & pix_x <=434 & pix_y >= 124 & pix_y <=124 ) | (pix_x >= 380 & pix_x <=435 & pix_y >= 125 & pix_y <=125 ) | (pix_x >= 382 & pix_x <=435 & pix_y >= 126 & pix_y <=126 ) | (pix_x >= 382 & pix_x <=436 & pix_y >= 127 & pix_y <=127 ) | (pix_x >= 382 & pix_x <=436 & pix_y >= 128 & pix_y <=128 ) | (pix_x >= 382 & pix_x <=437 & pix_y >= 129 & pix_y <=129 ) | (pix_x >= 382 & pix_x <=438 & pix_y >= 130 & pix_y <=130 ) | (pix_x >= 383 & pix_x <=440 & pix_y >= 131 & pix_y <=131 ) | (pix_x >= 385 & pix_x <=441 & pix_y >= 132 & pix_y <=132 ) | (pix_x >= 385 & pix_x <=442 & pix_y >= 133 & pix_y <=133 ) | (pix_x >= 385 & pix_x <=443 & pix_y >= 134 & pix_y <=134 ) | (pix_x >= 385 & pix_x <=445 & pix_y >= 135 & pix_y <=135 ) | (pix_x >= 383 & pix_x <=446 & pix_y >= 136 & pix_y <=136 ) | (pix_x >= 383 & pix_x <=446 & pix_y >= 137 & pix_y <=137 ) | (pix_x >= 383 & pix_x <=447 & pix_y >= 138 & pix_y <=138 ) | (pix_x >= 382 & pix_x <=448 & pix_y >= 139 & pix_y <=139 ) | (pix_x >= 382 & pix_x <=449 & pix_y >= 140 & pix_y <=140 ) | (pix_x >= 382 & pix_x <=383 & pix_y >= 141 & pix_y <=141 ) | (pix_x >= 385 & pix_x <=449 & pix_y >= 141 & pix_y <=141 ) | (pix_x >= 381 & pix_x <=383 & pix_y >= 142 & pix_y <=142 ) | (pix_x >= 385 & pix_x <=449 & pix_y >= 142 & pix_y <=142 ) | (pix_x >= 381 & pix_x <=383 & pix_y >= 143 & pix_y <=143 ) | (pix_x >= 385 & pix_x <=450 & pix_y >= 143 & pix_y <=143 ) | (pix_x >= 393 & pix_x <=450 & pix_y >= 144 & pix_y <=144 ) | (pix_x >= 393 & pix_x <=450 & pix_y >= 145 & pix_y <=145 ) | (pix_x >= 393 & pix_x <=451 & pix_y >= 146 & pix_y <=146 ) | (pix_x >= 393 & pix_x <=452 & pix_y >= 147 & pix_y <=147 ) | (pix_x >= 374 & pix_x <=376 & pix_y >= 148 & pix_y <=148 ) | (pix_x >= 393 & pix_x <=452 & pix_y >= 148 & pix_y <=148 ) | (pix_x >= 373 & pix_x <=375 & pix_y >= 149 & pix_y <=149 ) | (pix_x >= 393 & pix_x <=453 & pix_y >= 149 & pix_y <=149 ) | (pix_x >= 373 & pix_x <=374 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 393 & pix_x <=403 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 408 & pix_x <=454 & pix_y >= 150 & pix_y <=150 ) | (pix_x >= 393 & pix_x <=403 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 409 & pix_x <=454 & pix_y >= 151 & pix_y <=151 ) | (pix_x >= 385 & pix_x <=454 & pix_y >= 152 & pix_y <=151 ) | (pix_x >= 391 & pix_x <=395 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 401 & pix_x <=395 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 412 & pix_x <=454 & pix_y >= 152 & pix_y <=152 ) | (pix_x >= 387 & pix_x <=389 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 411 & pix_x <=455 & pix_y >= 153 & pix_y <=153 ) | (pix_x >= 387 & pix_x <=389 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 409 & pix_x <=413 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 417 & pix_x <=456 & pix_y >= 154 & pix_y <=154 ) | (pix_x >= 406 & pix_x <=411 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 417 & pix_x <=456 & pix_y >= 155 & pix_y <=155 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 415 & pix_x <=420 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 423 & pix_x <=457 & pix_y >= 156 & pix_y <=156 ) | (pix_x >= 414 & pix_x <=420 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 424 & pix_x <=457 & pix_y >= 157 & pix_y <=157 ) | (pix_x >= 411 & pix_x <=416 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 433 & pix_x <=457 & pix_y >= 158 & pix_y <=158 ) | (pix_x >= 409 & pix_x <=415 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 433 & pix_x <=458 & pix_y >= 159 & pix_y <=159 ) | (pix_x >= 407 & pix_x <=418 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 433 & pix_x <=458 & pix_y >= 160 & pix_y <=160 ) | (pix_x >= 407 & pix_x <=419 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 441 & pix_x <=458 & pix_y >= 161 & pix_y <=161 ) | (pix_x >= 407 & pix_x <=418 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 441 & pix_x <=458 & pix_y >= 162 & pix_y <=162 ) | (pix_x >= 405 & pix_x <=418 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 441 & pix_x <=418 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 443 & pix_x <=459 & pix_y >= 163 & pix_y <=163 ) | (pix_x >= 404 & pix_x <=420 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 444 & pix_x <=459 & pix_y >= 164 & pix_y <=164 ) | (pix_x >= 405 & pix_x <=421 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 165 & pix_y <=165 ) | (pix_x >= 409 & pix_x <=422 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 166 & pix_y <=166 ) | (pix_x >= 409 & pix_x <=429 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 445 & pix_x <=459 & pix_y >= 167 & pix_y <=167 ) | (pix_x >= 410 & pix_x <=435 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 445 & pix_x <=458 & pix_y >= 168 & pix_y <=168 ) | (pix_x >= 410 & pix_x <=440 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 446 & pix_x <=458 & pix_y >= 169 & pix_y <=169 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 436 & pix_x <=440 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 446 & pix_x <=459 & pix_y >= 170 & pix_y <=170 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 446 & pix_x <=458 & pix_y >= 171 & pix_y <=171 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 446 & pix_x <=458 & pix_y >= 172 & pix_y <=172 ) | (pix_x >= 410 & pix_x <=432 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 447 & pix_x <=456 & pix_y >= 173 & pix_y <=173 ) | (pix_x >= 411 & pix_x <=416 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 448 & pix_x <=456 & pix_y >= 174 & pix_y <=174 ) | (pix_x >= 412 & pix_x <=432 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 449 & pix_x <=456 & pix_y >= 175 & pix_y <=175 ) | (pix_x >= 414 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 444 & pix_x <=432 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 450 & pix_x <=455 & pix_y >= 176 & pix_y <=176 ) | (pix_x >= 414 & pix_x <=432 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 444 & pix_x <=445 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 451 & pix_x <=455 & pix_y >= 177 & pix_y <=177 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 422 & pix_x <=432 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 453 & pix_x <=455 & pix_y >= 178 & pix_y <=178 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 454 & pix_x <=446 & pix_y >= 179 & pix_y <=179 ) | (pix_x >= 374 & pix_x <=376 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 414 & pix_x <=416 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 423 & pix_x <=431 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 180 & pix_y <=180 ) | (pix_x >= 364 & pix_x <=376 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 415 & pix_x <=416 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 422 & pix_x <=431 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 181 & pix_y <=181 ) | (pix_x >= 356 & pix_x <=360 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 369 & pix_x <=376 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 422 & pix_x <=432 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 456 & pix_x <=457 & pix_y >= 182 & pix_y <=182 ) | (pix_x >= 353 & pix_x <=376 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 415 & pix_x <=418 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 443 & pix_x <=448 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 456 & pix_x <=458 & pix_y >= 183 & pix_y <=183 ) | (pix_x >= 357 & pix_x <=380 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 421 & pix_x <=432 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 184 & pix_y <=184 ) | (pix_x >= 356 & pix_x <=380 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 407 & pix_x <=408 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 422 & pix_x <=432 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 443 & pix_x <=447 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 456 & pix_x <=459 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 465 & pix_x <=467 & pix_y >= 185 & pix_y <=185 ) | (pix_x >= 356 & pix_x <=381 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 406 & pix_x <=408 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 457 & pix_x <=459 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 463 & pix_x <=469 & pix_y >= 186 & pix_y <=186 ) | (pix_x >= 356 & pix_x <=381 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 457 & pix_x <=458 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 463 & pix_x <=464 & pix_y >= 187 & pix_y <=187 ) | (pix_x >= 357 & pix_x <=382 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 404 & pix_x <=408 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 423 & pix_x <=432 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 188 & pix_y <=188 ) | (pix_x >= 359 & pix_x <=384 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 402 & pix_x <=408 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 415 & pix_x <=417 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 423 & pix_x <=417 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 189 & pix_y <=189 ) | (pix_x >= 361 & pix_x <=386 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 401 & pix_x <=408 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 416 & pix_x <=417 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 422 & pix_x <=417 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 190 & pix_y <=190 ) | (pix_x >= 361 & pix_x <=387 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 402 & pix_x <=408 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 416 & pix_x <=417 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 422 & pix_x <=417 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 454 & pix_x <=455 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 462 & pix_x <=466 & pix_y >= 191 & pix_y <=191 ) | (pix_x >= 365 & pix_x <=389 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 404 & pix_x <=408 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 416 & pix_x <=418 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 427 & pix_x <=431 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 442 & pix_x <=445 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 454 & pix_x <=456 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 192 & pix_y <=192 ) | (pix_x >= 365 & pix_x <=391 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 404 & pix_x <=408 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 416 & pix_x <=419 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 421 & pix_x <=419 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 426 & pix_x <=432 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 454 & pix_x <=457 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 193 & pix_y <=193 ) | (pix_x >= 366 & pix_x <=392 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 416 & pix_x <=422 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 425 & pix_x <=432 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 454 & pix_x <=458 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 194 & pix_y <=194 ) | (pix_x >= 367 & pix_x <=393 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 416 & pix_x <=421 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 425 & pix_x <=433 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 442 & pix_x <=444 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 454 & pix_x <=460 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 195 & pix_y <=195 ) | (pix_x >= 370 & pix_x <=395 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 405 & pix_x <=408 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 416 & pix_x <=434 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 454 & pix_x <=466 & pix_y >= 196 & pix_y <=196 ) | (pix_x >= 371 & pix_x <=408 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 416 & pix_x <=436 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 197 & pix_y <=197 ) | (pix_x >= 372 & pix_x <=408 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 416 & pix_x <=437 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 198 & pix_y <=198 ) | (pix_x >= 372 & pix_x <=408 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 416 & pix_x <=431 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 433 & pix_x <=437 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 445 & pix_x <=446 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 448 & pix_x <=446 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 199 & pix_y <=199 ) | (pix_x >= 373 & pix_x <=409 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 441 & pix_x <=446 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 453 & pix_x <=446 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 456 & pix_x <=466 & pix_y >= 200 & pix_y <=200 ) | (pix_x >= 373 & pix_x <=409 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 444 & pix_x <=446 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 453 & pix_x <=446 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 456 & pix_x <=467 & pix_y >= 201 & pix_y <=201 ) | (pix_x >= 373 & pix_x <=409 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 445 & pix_x <=442 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 452 & pix_x <=453 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 456 & pix_x <=468 & pix_y >= 202 & pix_y <=202 ) | (pix_x >= 374 & pix_x <=409 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 441 & pix_x <=443 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 452 & pix_x <=454 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 457 & pix_x <=469 & pix_y >= 203 & pix_y <=203 ) | (pix_x >= 375 & pix_x <=409 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 416 & pix_x <=438 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 452 & pix_x <=454 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 457 & pix_x <=470 & pix_y >= 204 & pix_y <=204 ) | (pix_x >= 375 & pix_x <=409 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 416 & pix_x <=439 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 441 & pix_x <=444 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 452 & pix_x <=453 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 461 & pix_x <=471 & pix_y >= 205 & pix_y <=205 ) | (pix_x >= 377 & pix_x <=409 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 442 & pix_x <=443 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 451 & pix_x <=453 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 461 & pix_x <=472 & pix_y >= 206 & pix_y <=206 ) | (pix_x >= 377 & pix_x <=409 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 451 & pix_x <=452 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 462 & pix_x <=472 & pix_y >= 207 & pix_y <=207 ) | (pix_x >= 379 & pix_x <=409 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 452 & pix_x <=453 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 459 & pix_x <=473 & pix_y >= 208 & pix_y <=208 ) | (pix_x >= 379 & pix_x <=409 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 452 & pix_x <=453 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 459 & pix_x <=474 & pix_y >= 209 & pix_y <=209 ) | (pix_x >= 379 & pix_x <=409 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 452 & pix_x <=439 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 458 & pix_x <=475 & pix_y >= 210 & pix_y <=210 ) | (pix_x >= 380 & pix_x <=410 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 452 & pix_x <=439 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 457 & pix_x <=476 & pix_y >= 211 & pix_y <=211 ) | (pix_x >= 381 & pix_x <=410 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 417 & pix_x <=439 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 451 & pix_x <=452 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 457 & pix_x <=459 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 465 & pix_x <=477 & pix_y >= 212 & pix_y <=212 ) | (pix_x >= 382 & pix_x <=411 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 418 & pix_x <=439 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 451 & pix_x <=452 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 457 & pix_x <=459 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 465 & pix_x <=478 & pix_y >= 213 & pix_y <=213 ) | (pix_x >= 382 & pix_x <=411 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 419 & pix_x <=439 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 456 & pix_x <=458 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 465 & pix_x <=479 & pix_y >= 214 & pix_y <=214 ) | (pix_x >= 268 & pix_x <=479 & pix_y >= 215 & pix_y <=214 ) | (pix_x >= 382 & pix_x <=411 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 420 & pix_x <=439 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 455 & pix_x <=458 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 465 & pix_x <=480 & pix_y >= 215 & pix_y <=215 ) | (pix_x >= 259 & pix_x <=480 & pix_y >= 216 & pix_y <=215 ) | (pix_x >= 269 & pix_x <=480 & pix_y >= 216 & pix_y <=215 ) | (pix_x >= 385 & pix_x <=413 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 421 & pix_x <=439 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 453 & pix_x <=459 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 468 & pix_x <=481 & pix_y >= 216 & pix_y <=216 ) | (pix_x >= 259 & pix_x <=481 & pix_y >= 217 & pix_y <=216 ) | (pix_x >= 269 & pix_x <=481 & pix_y >= 217 & pix_y <=216 ) | (pix_x >= 385 & pix_x <=414 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 423 & pix_x <=439 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 453 & pix_x <=459 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 468 & pix_x <=481 & pix_y >= 217 & pix_y <=217 ) | (pix_x >= 259 & pix_x <=481 & pix_y >= 218 & pix_y <=217 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 385 & pix_x <=416 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 425 & pix_x <=438 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 453 & pix_x <=461 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 468 & pix_x <=482 & pix_y >= 218 & pix_y <=218 ) | (pix_x >= 260 & pix_x <=482 & pix_y >= 219 & pix_y <=218 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 385 & pix_x <=418 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 427 & pix_x <=438 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 453 & pix_x <=466 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 468 & pix_x <=483 & pix_y >= 219 & pix_y <=219 ) | (pix_x >= 270 & pix_x <=483 & pix_y >= 220 & pix_y <=219 ) | (pix_x >= 387 & pix_x <=419 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 428 & pix_x <=439 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 453 & pix_x <=483 & pix_y >= 220 & pix_y <=220 ) | (pix_x >= 261 & pix_x <=483 & pix_y >= 221 & pix_y <=220 ) | (pix_x >= 387 & pix_x <=421 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 432 & pix_x <=439 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 448 & pix_x <=439 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 453 & pix_x <=484 & pix_y >= 221 & pix_y <=221 ) | (pix_x >= 261 & pix_x <=484 & pix_y >= 222 & pix_y <=221 ) | (pix_x >= 388 & pix_x <=424 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 453 & pix_x <=484 & pix_y >= 222 & pix_y <=222 ) | (pix_x >= 261 & pix_x <=262 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 273 & pix_x <=262 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 388 & pix_x <=429 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 453 & pix_x <=485 & pix_y >= 223 & pix_y <=223 ) | (pix_x >= 393 & pix_x <=431 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 224 & pix_y <=224 ) | (pix_x >= 393 & pix_x <=429 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 225 & pix_y <=225 ) | (pix_x >= 275 & pix_x <=276 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 395 & pix_x <=427 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 226 & pix_y <=226 ) | (pix_x >= 275 & pix_x <=276 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 397 & pix_x <=426 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 455 & pix_x <=485 & pix_y >= 227 & pix_y <=227 ) | (pix_x >= 265 & pix_x <=485 & pix_y >= 228 & pix_y <=227 ) | (pix_x >= 398 & pix_x <=400 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 403 & pix_x <=424 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 456 & pix_x <=485 & pix_y >= 228 & pix_y <=228 ) | (pix_x >= 265 & pix_x <=485 & pix_y >= 229 & pix_y <=228 ) | (pix_x >= 395 & pix_x <=425 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 429 & pix_x <=435 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 456 & pix_x <=472 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 474 & pix_x <=485 & pix_y >= 229 & pix_y <=229 ) | (pix_x >= 265 & pix_x <=266 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 393 & pix_x <=435 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 456 & pix_x <=470 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 475 & pix_x <=485 & pix_y >= 230 & pix_y <=230 ) | (pix_x >= 266 & pix_x <=268 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 393 & pix_x <=435 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 456 & pix_x <=469 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 476 & pix_x <=485 & pix_y >= 231 & pix_y <=231 ) | (pix_x >= 288 & pix_x <=289 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 399 & pix_x <=435 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 456 & pix_x <=464 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 477 & pix_x <=484 & pix_y >= 232 & pix_y <=232 ) | (pix_x >= 268 & pix_x <=269 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 289 & pix_x <=290 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 399 & pix_x <=435 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 457 & pix_x <=461 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 477 & pix_x <=484 & pix_y >= 233 & pix_y <=233 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 289 & pix_x <=292 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 458 & pix_x <=436 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 478 & pix_x <=484 & pix_y >= 234 & pix_y <=234 ) | (pix_x >= 269 & pix_x <=270 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 291 & pix_x <=293 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 481 & pix_x <=484 & pix_y >= 235 & pix_y <=235 ) | (pix_x >= 270 & pix_x <=484 & pix_y >= 236 & pix_y <=235 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 481 & pix_x <=483 & pix_y >= 236 & pix_y <=236 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 481 & pix_x <=483 & pix_y >= 237 & pix_y <=237 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 481 & pix_x <=482 & pix_y >= 238 & pix_y <=238 ) | (pix_x >= 280 & pix_x <=281 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 399 & pix_x <=436 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 481 & pix_x <=436 & pix_y >= 239 & pix_y <=239 ) | (pix_x >= 273 & pix_x <=436 & pix_y >= 240 & pix_y <=239 ) | (pix_x >= 279 & pix_x <=280 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 400 & pix_x <=437 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 481 & pix_x <=437 & pix_y >= 240 & pix_y <=240 ) | (pix_x >= 278 & pix_x <=280 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 401 & pix_x <=437 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 454 & pix_x <=459 & pix_y >= 241 & pix_y <=241 ) | (pix_x >= 277 & pix_x <=281 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 401 & pix_x <=438 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 454 & pix_x <=460 & pix_y >= 242 & pix_y <=242 ) | (pix_x >= 276 & pix_x <=282 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 401 & pix_x <=439 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 458 & pix_x <=460 & pix_y >= 243 & pix_y <=243 ) | (pix_x >= 277 & pix_x <=282 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 401 & pix_x <=442 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 457 & pix_x <=461 & pix_y >= 244 & pix_y <=244 ) | (pix_x >= 278 & pix_x <=282 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 401 & pix_x <=448 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 457 & pix_x <=462 & pix_y >= 245 & pix_y <=245 ) | (pix_x >= 279 & pix_x <=282 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 401 & pix_x <=462 & pix_y >= 246 & pix_y <=246 ) | (pix_x >= 279 & pix_x <=282 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 401 & pix_x <=464 & pix_y >= 247 & pix_y <=247 ) | (pix_x >= 399 & pix_x <=464 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 466 & pix_x <=467 & pix_y >= 248 & pix_y <=248 ) | (pix_x >= 399 & pix_x <=467 & pix_y >= 249 & pix_y <=249 ) | (pix_x >= 399 & pix_x <=466 & pix_y >= 250 & pix_y <=250 ) | (pix_x >= 399 & pix_x <=466 & pix_y >= 251 & pix_y <=251 ) | (pix_x >= 400 & pix_x <=466 & pix_y >= 252 & pix_y <=252 ) | (pix_x >= 400 & pix_x <=465 & pix_y >= 253 & pix_y <=253 ) | (pix_x >= 401 & pix_x <=465 & pix_y >= 254 & pix_y <=254 ) | (pix_x >= 402 & pix_x <=464 & pix_y >= 255 & pix_y <=255 ) | (pix_x >= 405 & pix_x <=465 & pix_y >= 256 & pix_y <=256 ) | (pix_x >= 405 & pix_x <=465 & pix_y >= 257 & pix_y <=257 ) | (pix_x >= 406 & pix_x <=432 & pix_y >= 258 & pix_y <=258 ) | (pix_x >= 439 & pix_x <=465 & pix_y >= 258 & pix_y <=258 ) | (pix_x >= 407 & pix_x <=416 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 418 & pix_x <=428 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 259 & pix_y <=259 ) | (pix_x >= 417 & pix_x <=420 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 260 & pix_y <=260 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 261 & pix_y <=261 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 262 & pix_y <=261 ) | (pix_x >= 444 & pix_x <=465 & pix_y >= 262 & pix_y <=262 ) | (pix_x >= 440 & pix_x <=465 & pix_y >= 263 & pix_y <=262 ) | (pix_x >= 444 & pix_x <=451 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 458 & pix_x <=465 & pix_y >= 263 & pix_y <=263 ) | (pix_x >= 409 & pix_x <=410 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 454 & pix_x <=457 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 460 & pix_x <=467 & pix_y >= 264 & pix_y <=264 ) | (pix_x >= 453 & pix_x <=458 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 461 & pix_x <=466 & pix_y >= 265 & pix_y <=265 ) | (pix_x >= 451 & pix_x <=459 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 463 & pix_x <=466 & pix_y >= 266 & pix_y <=266 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 463 & pix_x <=465 & pix_y >= 267 & pix_y <=267 ) | (pix_x >= 455 & pix_x <=460 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 463 & pix_x <=465 & pix_y >= 268 & pix_y <=268 ) | (pix_x >= 458 & pix_x <=464 & pix_y >= 269 & pix_y <=269 ) | (pix_x >= 457 & pix_x <=464 & pix_y >= 270 & pix_y <=269 ) | (pix_x >= 461 & pix_x <=464 & pix_y >= 270 & pix_y <=270 ) | (pix_x >= 457 & pix_x <=464 & pix_y >= 271 & pix_y <=270 ) | (pix_x >= 462 & pix_x <=464 & pix_y >= 271 & pix_y <=271 ) | (pix_x >= 432 & pix_x <=449 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 457 & pix_x <=449 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 461 & pix_x <=462 & pix_y >= 272 & pix_y <=272 ) | (pix_x >= 419 & pix_x <=423 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 433 & pix_x <=451 & pix_y >= 273 & pix_y <=273 ) | (pix_x >= 417 & pix_x <=429 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 438 & pix_x <=453 & pix_y >= 274 & pix_y <=274 ) | (pix_x >= 416 & pix_x <=423 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 425 & pix_x <=434 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 441 & pix_x <=456 & pix_y >= 275 & pix_y <=275 ) | (pix_x >= 415 & pix_x <=422 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 425 & pix_x <=436 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 441 & pix_x <=459 & pix_y >= 276 & pix_y <=276 ) | (pix_x >= 414 & pix_x <=428 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 430 & pix_x <=438 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 444 & pix_x <=460 & pix_y >= 277 & pix_y <=277 ) | (pix_x >= 413 & pix_x <=427 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 433 & pix_x <=440 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 446 & pix_x <=460 & pix_y >= 278 & pix_y <=278 ) | (pix_x >= 413 & pix_x <=422 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 435 & pix_x <=440 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 447 & pix_x <=459 & pix_y >= 279 & pix_y <=279 ) | (pix_x >= 412 & pix_x <=424 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 438 & pix_x <=441 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 449 & pix_x <=460 & pix_y >= 280 & pix_y <=280 ) | (pix_x >= 412 & pix_x <=424 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 439 & pix_x <=441 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 449 & pix_x <=459 & pix_y >= 281 & pix_y <=281 ) | (pix_x >= 412 & pix_x <=424 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 451 & pix_x <=459 & pix_y >= 282 & pix_y <=282 ) | (pix_x >= 412 & pix_x <=424 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 452 & pix_x <=458 & pix_y >= 283 & pix_y <=283 ) | (pix_x >= 413 & pix_x <=424 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 447 & pix_x <=457 & pix_y >= 284 & pix_y <=284 ) | (pix_x >= 417 & pix_x <=419 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 449 & pix_x <=456 & pix_y >= 285 & pix_y <=285 ) | (pix_x >= 456 & pix_x <=456 & pix_y >= 286 & pix_y <=285 ) | (pix_x >= 416 & pix_x <=419 & pix_y >= 288 & pix_y <=288 ) | (pix_x >= 429 & pix_x <=419 & pix_y >= 292 & pix_y <=288 ) | (pix_x >= 441 & pix_x <=442 & pix_y >= 292 & pix_y <=292 ) | (pix_x >= 427 & pix_x <=432 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 435 & pix_x <=444 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 449 & pix_x <=444 & pix_y >= 293 & pix_y <=293 ) | (pix_x >= 426 & pix_x <=445 & pix_y >= 294 & pix_y <=294 ) | (pix_x >= 447 & pix_x <=448 & pix_y >= 294 & pix_y <=294 ) | (pix_x >= 422 & pix_x <=424 & pix_y >= 295 & pix_y <=295 ) | (pix_x >= 426 & pix_x <=448 & pix_y >= 295 & pix_y <=295 ) | (pix_x >= 421 & pix_x <=448 & pix_y >= 296 & pix_y <=296 ) | (pix_x >= 421 & pix_x <=447 & pix_y >= 297 & pix_y <=297 ) | (pix_x >= 420 & pix_x <=447 & pix_y >= 298 & pix_y <=298 ) | (pix_x >= 420 & pix_x <=447 & pix_y >= 299 & pix_y <=299 ) | (pix_x >= 420 & pix_x <=447 & pix_y >= 300 & pix_y <=300 ) | (pix_x >= 420 & pix_x <=447 & pix_y >= 301 & pix_y <=301 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 302 & pix_y <=302 ) | (pix_x >= 420 & pix_x <=448 & pix_y >= 303 & pix_y <=303 ) | (pix_x >= 421 & pix_x <=448 & pix_y >= 304 & pix_y <=304 ) | (pix_x >= 421 & pix_x <=448 & pix_y >= 305 & pix_y <=305 ) | (pix_x >= 422 & pix_x <=448 & pix_y >= 306 & pix_y <=306 ) | (pix_x >= 423 & pix_x <=448 & pix_y >= 307 & pix_y <=307 ) | (pix_x >= 425 & pix_x <=448 & pix_y >= 308 & pix_y <=308 ) | (pix_x >= 425 & pix_x <=448 & pix_y >= 309 & pix_y <=309 ) | (pix_x >= 429 & pix_x <=442 & pix_y >= 310 & pix_y <=310 ) | (pix_x >= 444 & pix_x <=448 & pix_y >= 310 & pix_y <=310 ) | (pix_x >= 433 & pix_x <=442 & pix_y >= 311 & pix_y <=311 ) | (pix_x >= 445 & pix_x <=448 & pix_y >= 311 & pix_y <=311 ) | (pix_x >= 436 & pix_x <=437 & pix_y >= 312 & pix_y <=312 ) | (pix_x >= 445 & pix_x <=447 & pix_y >= 312 & pix_y <=312 ) | (pix_x >= 444 & pix_x <=446 & pix_y >= 313 & pix_y <=313 ) | (pix_x >= 444 & pix_x <=446 & pix_y >= 314 & pix_y <=314 ) | (pix_x >= 443 & pix_x <=446 & pix_y >= 315 & pix_y <=315 ) | (pix_x >= 443 & pix_x <=445 & pix_y >= 316 & pix_y <=316 ) | (pix_x >= 443 & pix_x <=444 & pix_y >= 317 & pix_y <=317 ) | (pix_x >= 348 & pix_x <=349 & pix_y >= 363 & pix_y <=363 ) | (pix_x >= 348 & pix_x <=349 & pix_y >= 364 & pix_y <=364 ) | (pix_x >= 348 & pix_x <=349 & pix_y >= 365 & pix_y <=365 ) | (pix_x >= 347 & pix_x <=349 & pix_y >= 368 & pix_y <=365 ) | (pix_x >= 346 & pix_x <=347 & pix_y >= 369 & pix_y <=369 ) | (pix_x >= 346 & pix_x <=347 & pix_y >= 370 & pix_y <=370 ) | (pix_x >= 345 & pix_x <=347 & pix_y >= 371 & pix_y <=370 ) | (pix_x >= 345 & pix_x <=347 & pix_y >= 372 & pix_y <=370 ) | (pix_x >= 341 & pix_x <=347 & pix_y >= 376 & pix_y <=370 ) | (pix_x >= 339 & pix_x <=347 & pix_y >= 380 & pix_y <=370 ) | (pix_x >= 337 & pix_x <=347 & pix_y >= 383 & pix_y <=370 ) | (pix_x >= 333 & pix_x <=347 & pix_y >= 391 & pix_y <=370 ) | (pix_x >= 272 & pix_x <=347 & pix_y >= 392 & pix_y <=370 ) | (pix_x >= 332 & pix_x <=333 & pix_y >= 392 & pix_y <=392 ) | (pix_x >= 272 & pix_x <=333 & pix_y >= 393 & pix_y <=392 ) | (pix_x >= 332 & pix_x <=333 & pix_y >= 393 & pix_y <=392 ) | (pix_x >= 272 & pix_x <=333 & pix_y >= 394 & pix_y <=392 ) | (pix_x >= 332 & pix_x <=333 & pix_y >= 394 & pix_y <=392 ) | (pix_x >= 329 & pix_x <=330 & pix_y >= 395 & pix_y <=395 ) | (pix_x >= 275 & pix_x <=330 & pix_y >= 396 & pix_y <=395 ) | (pix_x >= 329 & pix_x <=331 & pix_y >= 396 & pix_y <=396 ) | (pix_x >= 275 & pix_x <=276 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 326 & pix_x <=328 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 330 & pix_x <=331 & pix_y >= 397 & pix_y <=397 ) | (pix_x >= 275 & pix_x <=277 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 280 & pix_x <=277 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 324 & pix_x <=328 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 330 & pix_x <=328 & pix_y >= 398 & pix_y <=398 ) | (pix_x >= 275 & pix_x <=277 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 280 & pix_x <=277 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 323 & pix_x <=328 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 330 & pix_x <=328 & pix_y >= 399 & pix_y <=399 ) | (pix_x >= 275 & pix_x <=279 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 281 & pix_x <=282 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 287 & pix_x <=300 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 321 & pix_x <=330 & pix_y >= 400 & pix_y <=400 ) | (pix_x >= 275 & pix_x <=279 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 281 & pix_x <=283 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 286 & pix_x <=301 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 321 & pix_x <=330 & pix_y >= 401 & pix_y <=401 ) | (pix_x >= 275 & pix_x <=279 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 281 & pix_x <=302 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 316 & pix_x <=329 & pix_y >= 402 & pix_y <=402 ) | (pix_x >= 276 & pix_x <=304 & pix_y >= 403 & pix_y <=403 ) | (pix_x >= 313 & pix_x <=329 & pix_y >= 403 & pix_y <=403 ) | (pix_x >= 277 & pix_x <=329 & pix_y >= 404 & pix_y <=404 ) | (pix_x >= 277 & pix_x <=328 & pix_y >= 405 & pix_y <=405 ) | (pix_x >= 277 & pix_x <=328 & pix_y >= 406 & pix_y <=406 ) | (pix_x >= 277 & pix_x <=328 & pix_y >= 407 & pix_y <=407 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 408 & pix_y <=408 ) | (pix_x >= 278 & pix_x <=328 & pix_y >= 409 & pix_y <=409 ) | (pix_x >= 279 & pix_x <=327 & pix_y >= 410 & pix_y <=410 ) | (pix_x >= 279 & pix_x <=327 & pix_y >= 411 & pix_y <=411 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 412 & pix_y <=412 ) | (pix_x >= 280 & pix_x <=327 & pix_y >= 413 & pix_y <=413 ) | (pix_x >= 426 & pix_x <=428 & pix_y >= 413 & pix_y <=413 ) | (pix_x >= 281 & pix_x <=326 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 414 & pix_y <=414 ) | (pix_x >= 281 & pix_x <=326 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 415 & pix_y <=415 ) | (pix_x >= 281 & pix_x <=326 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 416 & pix_y <=416 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 417 & pix_y <=417 ) | (pix_x >= 282 & pix_x <=326 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 426 & pix_x <=429 & pix_y >= 418 & pix_y <=418 ) | (pix_x >= 283 & pix_x <=326 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 427 & pix_x <=429 & pix_y >= 419 & pix_y <=419 ) | (pix_x >= 283 & pix_x <=325 & pix_y >= 420 & pix_y <=420 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 426 & pix_x <=427 & pix_y >= 421 & pix_y <=421 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 422 & pix_y <=422 ) | (pix_x >= 284 & pix_x <=325 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 425 & pix_x <=429 & pix_y >= 423 & pix_y <=423 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 424 & pix_y <=424 ) | (pix_x >= 285 & pix_x <=324 & pix_y >= 425 & pix_y <=425 ) | (pix_x >= 286 & pix_x <=323 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 425 & pix_x <=426 & pix_y >= 426 & pix_y <=426 ) | (pix_x >= 286 & pix_x <=322 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 427 & pix_y <=427 ) | (pix_x >= 287 & pix_x <=322 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 425 & pix_x <=427 & pix_y >= 428 & pix_y <=428 ) | (pix_x >= 288 & pix_x <=321 & pix_y >= 429 & pix_y <=429 ) | (pix_x >= 288 & pix_x <=321 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 424 & pix_x <=425 & pix_y >= 430 & pix_y <=430 ) | (pix_x >= 288 & pix_x <=320 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 424 & pix_x <=426 & pix_y >= 431 & pix_y <=431 ) | (pix_x >= 289 & pix_x <=319 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 425 & pix_x <=428 & pix_y >= 432 & pix_y <=432 ) | (pix_x >= 289 & pix_x <=319 & pix_y >= 433 & pix_y <=433 ) | (pix_x >= 290 & pix_x <=318 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 424 & pix_x <=318 & pix_y >= 434 & pix_y <=434 ) | (pix_x >= 291 & pix_x <=318 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 423 & pix_x <=425 & pix_y >= 435 & pix_y <=435 ) | (pix_x >= 291 & pix_x <=317 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 424 & pix_x <=426 & pix_y >= 436 & pix_y <=436 ) | (pix_x >= 292 & pix_x <=316 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 425 & pix_x <=316 & pix_y >= 437 & pix_y <=437 ) | (pix_x >= 292 & pix_x <=315 & pix_y >= 438 & pix_y <=438 ) | (pix_x >= 292 & pix_x <=314 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 439 & pix_y <=439 ) | (pix_x >= 293 & pix_x <=313 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 423 & pix_x <=425 & pix_y >= 440 & pix_y <=440 ) | (pix_x >= 293 & pix_x <=313 & pix_y >= 441 & pix_y <=441 ) | (pix_x >= 294 & pix_x <=312 & pix_y >= 442 & pix_y <=442 ) | (pix_x >= 294 & pix_x <=311 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 422 & pix_x <=423 & pix_y >= 443 & pix_y <=443 ) | (pix_x >= 295 & pix_x <=310 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 422 & pix_x <=423 & pix_y >= 444 & pix_y <=444 ) | (pix_x >= 295 & pix_x <=310 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 423 & pix_x <=424 & pix_y >= 445 & pix_y <=445 ) | (pix_x >= 296 & pix_x <=309 & pix_y >= 446 & pix_y <=446 ) | (pix_x >= 296 & pix_x <=309 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 421 & pix_x <=309 & pix_y >= 447 & pix_y <=447 ) | (pix_x >= 297 & pix_x <=298 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 300 & pix_x <=308 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 421 & pix_x <=422 & pix_y >= 448 & pix_y <=448 ) | (pix_x >= 300 & pix_x <=308 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 421 & pix_x <=424 & pix_y >= 449 & pix_y <=449 ) | (pix_x >= 299 & pix_x <=307 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 424 & pix_x <=307 & pix_y >= 450 & pix_y <=450 ) | (pix_x >= 300 & pix_x <=306 & pix_y >= 451 & pix_y <=451 ) | (pix_x >= 300 & pix_x <=301 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 304 & pix_x <=306 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 420 & pix_x <=422 & pix_y >= 452 & pix_y <=452 ) | (pix_x >= 301 & pix_x <=305 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 420 & pix_x <=423 & pix_y >= 453 & pix_y <=453 ) | (pix_x >= 302 & pix_x <=303 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 421 & pix_x <=423 & pix_y >= 454 & pix_y <=454 ) | (pix_x >= 302 & pix_x <=303 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 420 & pix_x <=303 & pix_y >= 455 & pix_y <=455 ) | (pix_x >= 303 & pix_x <=304 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=421 & pix_y >= 456 & pix_y <=456 ) | (pix_x >= 304 & pix_x <=421 & pix_y >= 457 & pix_y <=456 ) | (pix_x >= 419 & pix_x <=422 & pix_y >= 457 & pix_y <=457 ) | (pix_x >= 420 & pix_x <=423 & pix_y >= 458 & pix_y <=458 ) | (pix_x >= 418 & pix_x <=420 & pix_y >= 461 & pix_y <=461 ) | (pix_x >= 419 & pix_x <=420 & pix_y >= 462 & pix_y <=462 ) ;



endmodule
