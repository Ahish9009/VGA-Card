module pixel_itr(
    input wire clk,
    input wire pix_clk,
    input wire rst,
    output wire [9:0] pix_x,
    output wire [9:0] pix_y,
    output wire h_sync,
    output wire v_sync,
    output wire draw_active,
    output wire screen_end,
    output wire draw_end
    );
	 
	// FOR 800 X 600
    // parameter h_sync_strt = 56;          
    // parameter h_sync_end  = 56 + 120;         
    // parameter v_sync_strt = 600 + 37;        
    // parameter v_sync_end  = 600 + 37 + 6;   
    // parameter h_draw_min  = 56 + 120 + 64;   
    // parameter v_draw_max  = 600 - 1;            
    // parameter h_max = 1040;           
    // parameter v_max = 666 - 1;
	 
	// FOR 640 X 480
    parameter h_sync_strt = 16;          
    parameter h_sync_end  = 16 + 96;         
    parameter v_sync_strt = 480 + 10;        
    parameter v_sync_end  = 480 + 10 + 2;   
    parameter h_draw_min  = 16 + 96 + 48;   
    parameter v_draw_max  = 480 - 1;            
    parameter h_max = 800;           
    parameter v_max = 525 - 1;

    reg [9:0] h_pos=0;
	 reg [9:0] v_pos=0; 
	
    // --------------- SYNC SIGNALS BLOCK ---------------
    assign h_sync = (h_pos >= h_sync_strt && h_pos < h_sync_end) ? 0 : 1;
    assign v_sync = (v_pos >= v_sync_strt && v_pos < v_sync_end) ? 0 : 1;
    // --------------------------------------------------
		
	// -------------- PIXEL POSITION BLOCK --------------
    // assign pix_x = (h_pos >= h_draw_min) ? h_pos : 0;        
    assign pix_x = (h_pos >= h_draw_min) ? h_pos - h_draw_min : 0;        
	 assign pix_y = (v_pos <= v_draw_max) ? v_pos : v_draw_max;        
    // --------------------------------------------------

    // -------- BLANKING / DRAWING PERIOD BLOCK ---------
    assign draw_active = (h_pos < h_draw_min | v_pos > v_draw_max) ? 0 : 1;
    // --------------------------------------------------

    // ----------------- LIMITS BLOCK -------------------
    assign screen_end = (h_pos == h_max & v_pos == v_max);
    assign draw_end = (h_pos == h_max & v_pos == v_draw_max);
    // --------------------------------------------------
    
    // ------------------ MAIN BLOCK --------------------
    always @ (posedge clk) begin
        if (rst) begin
            h_pos <= 0; 
            v_pos <= 0;
        end

        if(pix_clk) begin
            if (h_pos < h_max) begin
                h_pos <= h_pos + 1; 
            end
            else begin
                h_pos <= 0;
                v_pos <= v_pos + 1;
            end

            if (v_pos == v_max) begin
                    v_pos <= 0;
            end
        end
    end
    // --------------------------------------------------

endmodule

//////////////////////////////////////////////////////////////////////////////////

module screen_design(
	input clk,
	input rst,
	output h_sync,
	output v_sync,
	output r_out,
	output g_out,
	output b_out
);

//---------------GENERATING PIXEL CLOCK----------------------
reg count = 0, pix_clk = 0;

always @(posedge clk) begin
	
	if (rst == 1) begin
		count <= 0;
		pix_clk <= 0;
	end 
	if (count == 1) begin
		pix_clk <= 1;
		count <= 0;
	end 
	else begin
		pix_clk <= 0;
		count <= count + 1;

	end
end

//-----------------------------------------------------------

//-------------GETTING CURRENT PIXEL COORDINATES-------------
wire [9:0] pix_x;
wire [9:0] pix_y;

pixel_itr show(
	.clk(clk),
   .pix_clk(pix_clk),
	.rst(rst),
	.pix_x(pix_x),
	.pix_y(pix_y),
	.h_sync(h_sync),
	.v_sync(v_sync)
);
//-----------------------------------------------------------

//----------GENERATING WINDOWS LOGO(4 SQUARES)---------------

wire win1, win2, win3, win4;
assign win1 = (pix_x == 17 & pix_y == 297)| (pix_x == 17 & pix_y == 298)| (pix_x == 18 & pix_y == 297)| (pix_x == 18 & pix_y == 298)| (pix_x == 19 & pix_y == 297)| (pix_x == 19 & pix_y == 298)| (pix_x == 19 & pix_y == 299)| (pix_x == 19 & pix_y == 300)| (pix_x == 19 & pix_y == 301)| (pix_x == 19 & pix_y == 302)| (pix_x == 19 & pix_y == 303)| (pix_x == 19 & pix_y == 304)| (pix_x == 19 & pix_y == 323)| (pix_x == 19 & pix_y == 324)| (pix_x == 19 & pix_y == 325)| (pix_x == 19 & pix_y == 326)| (pix_x == 20 & pix_y == 297)| (pix_x == 20 & pix_y == 298)| (pix_x == 20 & pix_y == 299)| (pix_x == 20 & pix_y == 300)| (pix_x == 20 & pix_y == 301)| (pix_x == 20 & pix_y == 302)| (pix_x == 20 & pix_y == 303)| (pix_x == 20 & pix_y == 304)| (pix_x == 20 & pix_y == 323)| (pix_x == 20 & pix_y == 324)| (pix_x == 20 & pix_y == 325)| (pix_x == 20 & pix_y == 326)| (pix_x == 21 & pix_y == 297)| (pix_x == 21 & pix_y == 298)| (pix_x == 21 & pix_y == 299)| (pix_x == 21 & pix_y == 300)| (pix_x == 21 & pix_y == 301)| (pix_x == 21 & pix_y == 302)| (pix_x == 21 & pix_y == 303)| (pix_x == 21 & pix_y == 304)| (pix_x == 21 & pix_y == 323)| (pix_x == 21 & pix_y == 324)| (pix_x == 21 & pix_y == 325)| (pix_x == 21 & pix_y == 326)| (pix_x == 22 & pix_y == 297)| (pix_x == 22 & pix_y == 298)| (pix_x == 22 & pix_y == 299)| (pix_x == 22 & pix_y == 300)| (pix_x == 22 & pix_y == 301)| (pix_x == 22 & pix_y == 302)| (pix_x == 22 & pix_y == 303)| (pix_x == 22 & pix_y == 304)| (pix_x == 22 & pix_y == 312)| (pix_x == 22 & pix_y == 315)| (pix_x == 22 & pix_y == 316)| (pix_x == 22 & pix_y == 318)| (pix_x == 22 & pix_y == 319)| (pix_x == 22 & pix_y == 323)| (pix_x == 22 & pix_y == 324)| (pix_x == 22 & pix_y == 325)| (pix_x == 22 & pix_y == 326)| (pix_x == 22 & pix_y == 328)| (pix_x == 22 & pix_y == 329)| (pix_x == 23 & pix_y == 297)| (pix_x == 23 & pix_y == 298)| (pix_x == 23 & pix_y == 299)| (pix_x == 23 & pix_y == 300)| (pix_x == 23 & pix_y == 301)| (pix_x == 23 & pix_y == 302)| (pix_x == 23 & pix_y == 303)| (pix_x == 23 & pix_y == 304)| (pix_x == 23 & pix_y == 312)| (pix_x == 23 & pix_y == 315)| (pix_x == 23 & pix_y == 316)| (pix_x == 23 & pix_y == 318)| (pix_x == 23 & pix_y == 319)| (pix_x == 23 & pix_y == 323)| (pix_x == 23 & pix_y == 324)| (pix_x == 23 & pix_y == 325)| (pix_x == 23 & pix_y == 326)| (pix_x == 23 & pix_y == 328)| (pix_x == 23 & pix_y == 329)| (pix_x == 24 & pix_y == 290)| (pix_x == 24 & pix_y == 291)| (pix_x == 24 & pix_y == 297)| (pix_x == 24 & pix_y == 298)| (pix_x == 24 & pix_y == 299)| (pix_x == 24 & pix_y == 300)| (pix_x == 24 & pix_y == 301)| (pix_x == 24 & pix_y == 302)| (pix_x == 24 & pix_y == 303)| (pix_x == 24 & pix_y == 307)| (pix_x == 24 & pix_y == 310)| (pix_x == 24 & pix_y == 311)| (pix_x == 24 & pix_y == 312)| (pix_x == 24 & pix_y == 315)| (pix_x == 24 & pix_y == 316)| (pix_x == 24 & pix_y == 318)| (pix_x == 24 & pix_y == 319)| (pix_x == 24 & pix_y == 325)| (pix_x == 24 & pix_y == 326)| (pix_x == 24 & pix_y == 328)| (pix_x == 24 & pix_y == 329)| (pix_x == 25 & pix_y == 290)| (pix_x == 25 & pix_y == 291)| (pix_x == 25 & pix_y == 297)| (pix_x == 25 & pix_y == 298)| (pix_x == 25 & pix_y == 299)| (pix_x == 25 & pix_y == 300)| (pix_x == 25 & pix_y == 301)| (pix_x == 25 & pix_y == 302)| (pix_x == 25 & pix_y == 303)| (pix_x == 25 & pix_y == 307)| (pix_x == 25 & pix_y == 310)| (pix_x == 25 & pix_y == 311)| (pix_x == 25 & pix_y == 312)| (pix_x == 25 & pix_y == 315)| (pix_x == 25 & pix_y == 316)| (pix_x == 25 & pix_y == 318)| (pix_x == 25 & pix_y == 319)| (pix_x == 25 & pix_y == 325)| (pix_x == 25 & pix_y == 326)| (pix_x == 25 & pix_y == 328)| (pix_x == 25 & pix_y == 329)| (pix_x == 26 & pix_y == 290)| (pix_x == 26 & pix_y == 291)| (pix_x == 26 & pix_y == 299)| (pix_x == 26 & pix_y == 300)| (pix_x == 26 & pix_y == 301)| (pix_x == 26 & pix_y == 302)| (pix_x == 26 & pix_y == 303)| (pix_x == 26 & pix_y == 304)| (pix_x == 26 & pix_y == 307)| (pix_x == 26 & pix_y == 312)| (pix_x == 26 & pix_y == 313)| (pix_x == 26 & pix_y == 314)| (pix_x == 26 & pix_y == 315)| (pix_x == 26 & pix_y == 316)| (pix_x == 26 & pix_y == 318)| (pix_x == 26 & pix_y == 319)| (pix_x == 26 & pix_y == 323)| (pix_x == 26 & pix_y == 324)| (pix_x == 26 & pix_y == 325)| (pix_x == 26 & pix_y == 326)| (pix_x == 26 & pix_y == 332)| (pix_x == 26 & pix_y == 333)| (pix_x == 26 & pix_y == 334)| (pix_x == 26 & pix_y == 340)| (pix_x == 27 & pix_y == 290)| (pix_x == 27 & pix_y == 291)| (pix_x == 27 & pix_y == 299)| (pix_x == 27 & pix_y == 300)| (pix_x == 27 & pix_y == 301)| (pix_x == 27 & pix_y == 302)| (pix_x == 27 & pix_y == 303)| (pix_x == 27 & pix_y == 304)| (pix_x == 27 & pix_y == 307)| (pix_x == 27 & pix_y == 312)| (pix_x == 27 & pix_y == 313)| (pix_x == 27 & pix_y == 314)| (pix_x == 27 & pix_y == 315)| (pix_x == 27 & pix_y == 316)| (pix_x == 27 & pix_y == 318)| (pix_x == 27 & pix_y == 319)| (pix_x == 27 & pix_y == 323)| (pix_x == 27 & pix_y == 324)| (pix_x == 27 & pix_y == 325)| (pix_x == 27 & pix_y == 326)| (pix_x == 27 & pix_y == 332)| (pix_x == 27 & pix_y == 333)| (pix_x == 27 & pix_y == 334)| (pix_x == 27 & pix_y == 340)| (pix_x == 28 & pix_y == 290)| (pix_x == 28 & pix_y == 291)| (pix_x == 28 & pix_y == 299)| (pix_x == 28 & pix_y == 300)| (pix_x == 28 & pix_y == 301)| (pix_x == 28 & pix_y == 302)| (pix_x == 28 & pix_y == 303)| (pix_x == 28 & pix_y == 304)| (pix_x == 28 & pix_y == 307)| (pix_x == 28 & pix_y == 312)| (pix_x == 28 & pix_y == 313)| (pix_x == 28 & pix_y == 314)| (pix_x == 28 & pix_y == 315)| (pix_x == 28 & pix_y == 316)| (pix_x == 28 & pix_y == 318)| (pix_x == 28 & pix_y == 319)| (pix_x == 28 & pix_y == 323)| (pix_x == 28 & pix_y == 324)| (pix_x == 28 & pix_y == 325)| (pix_x == 28 & pix_y == 326)| (pix_x == 28 & pix_y == 332)| (pix_x == 28 & pix_y == 333)| (pix_x == 28 & pix_y == 334)| (pix_x == 28 & pix_y == 340)| (pix_x == 29 & pix_y == 289)| (pix_x == 29 & pix_y == 305)| (pix_x == 29 & pix_y == 306)| (pix_x == 29 & pix_y == 307)| (pix_x == 29 & pix_y == 308)| (pix_x == 29 & pix_y == 309)| (pix_x == 29 & pix_y == 318)| (pix_x == 29 & pix_y == 319)| (pix_x == 29 & pix_y == 320)| (pix_x == 29 & pix_y == 321)| (pix_x == 29 & pix_y == 333)| (pix_x == 29 & pix_y == 334)| (pix_x == 30 & pix_y == 289)| (pix_x == 30 & pix_y == 305)| (pix_x == 30 & pix_y == 306)| (pix_x == 30 & pix_y == 307)| (pix_x == 30 & pix_y == 308)| (pix_x == 30 & pix_y == 309)| (pix_x == 30 & pix_y == 318)| (pix_x == 30 & pix_y == 319)| (pix_x == 30 & pix_y == 320)| (pix_x == 30 & pix_y == 321)| (pix_x == 30 & pix_y == 333)| (pix_x == 30 & pix_y == 334)| (pix_x == 31 & pix_y == 289)| (pix_x == 31 & pix_y == 343)| (pix_x == 31 & pix_y == 344)| (pix_x == 32 & pix_y == 289)| (pix_x == 32 & pix_y == 343)| (pix_x == 32 & pix_y == 344)| (pix_x == 33 & pix_y == 289)| (pix_x == 33 & pix_y == 343)| (pix_x == 33 & pix_y == 344)| (pix_x == 34 & pix_y == 287)| (pix_x == 34 & pix_y == 288)| (pix_x == 34 & pix_y == 289)| (pix_x == 34 & pix_y == 294)| (pix_x == 34 & pix_y == 327)| (pix_x == 34 & pix_y == 341)| (pix_x == 34 & pix_y == 342)| (pix_x == 34 & pix_y == 343)| (pix_x == 34 & pix_y == 344)| (pix_x == 34 & pix_y == 345)| (pix_x == 34 & pix_y == 346)| (pix_x == 34 & pix_y == 347)| (pix_x == 34 & pix_y == 348)| (pix_x == 34 & pix_y == 349)| (pix_x == 34 & pix_y == 353)| (pix_x == 34 & pix_y == 354)| (pix_x == 35 & pix_y == 287)| (pix_x == 35 & pix_y == 288)| (pix_x == 35 & pix_y == 289)| (pix_x == 35 & pix_y == 294)| (pix_x == 35 & pix_y == 327)| (pix_x == 35 & pix_y == 341)| (pix_x == 35 & pix_y == 342)| (pix_x == 35 & pix_y == 343)| (pix_x == 35 & pix_y == 344)| (pix_x == 35 & pix_y == 345)| (pix_x == 35 & pix_y == 346)| (pix_x == 35 & pix_y == 347)| (pix_x == 35 & pix_y == 348)| (pix_x == 35 & pix_y == 349)| (pix_x == 35 & pix_y == 353)| (pix_x == 35 & pix_y == 354)| (pix_x == 36 & pix_y == 325)| (pix_x == 36 & pix_y == 326)| (pix_x == 36 & pix_y == 327)| (pix_x == 36 & pix_y == 328)| (pix_x == 36 & pix_y == 329)| (pix_x == 36 & pix_y == 336)| (pix_x == 36 & pix_y == 337)| (pix_x == 36 & pix_y == 340)| (pix_x == 36 & pix_y == 343)| (pix_x == 36 & pix_y == 344)| (pix_x == 36 & pix_y == 345)| (pix_x == 36 & pix_y == 346)| (pix_x == 36 & pix_y == 347)| (pix_x == 36 & pix_y == 348)| (pix_x == 36 & pix_y == 349)| (pix_x == 36 & pix_y == 350)| (pix_x == 36 & pix_y == 351)| (pix_x == 36 & pix_y == 352)| (pix_x == 36 & pix_y == 353)| (pix_x == 36 & pix_y == 354)| (pix_x == 36 & pix_y == 355)| (pix_x == 37 & pix_y == 325)| (pix_x == 37 & pix_y == 326)| (pix_x == 37 & pix_y == 327)| (pix_x == 37 & pix_y == 328)| (pix_x == 37 & pix_y == 329)| (pix_x == 37 & pix_y == 336)| (pix_x == 37 & pix_y == 337)| (pix_x == 37 & pix_y == 340)| (pix_x == 37 & pix_y == 343)| (pix_x == 37 & pix_y == 344)| (pix_x == 37 & pix_y == 345)| (pix_x == 37 & pix_y == 346)| (pix_x == 37 & pix_y == 347)| (pix_x == 37 & pix_y == 348)| (pix_x == 37 & pix_y == 349)| (pix_x == 37 & pix_y == 350)| (pix_x == 37 & pix_y == 351)| (pix_x == 37 & pix_y == 352)| (pix_x == 37 & pix_y == 353)| (pix_x == 37 & pix_y == 354)| (pix_x == 37 & pix_y == 355)| (pix_x == 38 & pix_y == 279)| (pix_x == 38 & pix_y == 280)| (pix_x == 38 & pix_y == 281)| (pix_x == 38 & pix_y == 320)| (pix_x == 38 & pix_y == 321)| (pix_x == 38 & pix_y == 327)| (pix_x == 38 & pix_y == 328)| (pix_x == 38 & pix_y == 329)| (pix_x == 38 & pix_y == 336)| (pix_x == 38 & pix_y == 337)| (pix_x == 38 & pix_y == 338)| (pix_x == 38 & pix_y == 339)| (pix_x == 38 & pix_y == 345)| (pix_x == 38 & pix_y == 346)| (pix_x == 38 & pix_y == 347)| (pix_x == 38 & pix_y == 348)| (pix_x == 38 & pix_y == 349)| (pix_x == 38 & pix_y == 350)| (pix_x == 38 & pix_y == 351)| (pix_x == 38 & pix_y == 352)| (pix_x == 38 & pix_y == 353)| (pix_x == 38 & pix_y == 354)| (pix_x == 38 & pix_y == 361)| (pix_x == 38 & pix_y == 362)| (pix_x == 39 & pix_y == 279)| (pix_x == 39 & pix_y == 280)| (pix_x == 39 & pix_y == 281)| (pix_x == 39 & pix_y == 320)| (pix_x == 39 & pix_y == 321)| (pix_x == 39 & pix_y == 327)| (pix_x == 39 & pix_y == 328)| (pix_x == 39 & pix_y == 329)| (pix_x == 39 & pix_y == 336)| (pix_x == 39 & pix_y == 337)| (pix_x == 39 & pix_y == 338)| (pix_x == 39 & pix_y == 339)| (pix_x == 39 & pix_y == 345)| (pix_x == 39 & pix_y == 346)| (pix_x == 39 & pix_y == 347)| (pix_x == 39 & pix_y == 348)| (pix_x == 39 & pix_y == 349)| (pix_x == 39 & pix_y == 350)| (pix_x == 39 & pix_y == 351)| (pix_x == 39 & pix_y == 352)| (pix_x == 39 & pix_y == 353)| (pix_x == 39 & pix_y == 354)| (pix_x == 39 & pix_y == 361)| (pix_x == 39 & pix_y == 362)| (pix_x == 40 & pix_y == 279)| (pix_x == 40 & pix_y == 280)| (pix_x == 40 & pix_y == 281)| (pix_x == 40 & pix_y == 320)| (pix_x == 40 & pix_y == 321)| (pix_x == 40 & pix_y == 327)| (pix_x == 40 & pix_y == 328)| (pix_x == 40 & pix_y == 329)| (pix_x == 40 & pix_y == 336)| (pix_x == 40 & pix_y == 337)| (pix_x == 40 & pix_y == 338)| (pix_x == 40 & pix_y == 339)| (pix_x == 40 & pix_y == 345)| (pix_x == 40 & pix_y == 346)| (pix_x == 40 & pix_y == 347)| (pix_x == 40 & pix_y == 348)| (pix_x == 40 & pix_y == 349)| (pix_x == 40 & pix_y == 350)| (pix_x == 40 & pix_y == 351)| (pix_x == 40 & pix_y == 352)| (pix_x == 40 & pix_y == 353)| (pix_x == 40 & pix_y == 354)| (pix_x == 40 & pix_y == 361)| (pix_x == 40 & pix_y == 362)| (pix_x == 41 & pix_y == 254)| (pix_x == 41 & pix_y == 255)| (pix_x == 41 & pix_y == 256)| (pix_x == 41 & pix_y == 353)| (pix_x == 41 & pix_y == 354)| (pix_x == 41 & pix_y == 355)| (pix_x == 41 & pix_y == 361)| (pix_x == 41 & pix_y == 362)| (pix_x == 41 & pix_y == 363)| (pix_x == 41 & pix_y == 364)| (pix_x == 42 & pix_y == 254)| (pix_x == 42 & pix_y == 255)| (pix_x == 42 & pix_y == 256)| (pix_x == 42 & pix_y == 353)| (pix_x == 42 & pix_y == 354)| (pix_x == 42 & pix_y == 355)| (pix_x == 42 & pix_y == 361)| (pix_x == 42 & pix_y == 362)| (pix_x == 42 & pix_y == 363)| (pix_x == 42 & pix_y == 364)| (pix_x == 43 & pix_y == 252)| (pix_x == 43 & pix_y == 253)| (pix_x == 43 & pix_y == 254)| (pix_x == 43 & pix_y == 255)| (pix_x == 43 & pix_y == 269)| (pix_x == 43 & pix_y == 270)| (pix_x == 43 & pix_y == 271)| (pix_x == 43 & pix_y == 272)| (pix_x == 43 & pix_y == 273)| (pix_x == 43 & pix_y == 294)| (pix_x == 43 & pix_y == 302)| (pix_x == 43 & pix_y == 303)| (pix_x == 43 & pix_y == 360)| (pix_x == 43 & pix_y == 361)| (pix_x == 43 & pix_y == 362)| (pix_x == 44 & pix_y == 252)| (pix_x == 44 & pix_y == 253)| (pix_x == 44 & pix_y == 254)| (pix_x == 44 & pix_y == 255)| (pix_x == 44 & pix_y == 269)| (pix_x == 44 & pix_y == 270)| (pix_x == 44 & pix_y == 271)| (pix_x == 44 & pix_y == 272)| (pix_x == 44 & pix_y == 273)| (pix_x == 44 & pix_y == 294)| (pix_x == 44 & pix_y == 302)| (pix_x == 44 & pix_y == 303)| (pix_x == 44 & pix_y == 360)| (pix_x == 44 & pix_y == 361)| (pix_x == 44 & pix_y == 362)| (pix_x == 45 & pix_y == 252)| (pix_x == 45 & pix_y == 253)| (pix_x == 45 & pix_y == 254)| (pix_x == 45 & pix_y == 255)| (pix_x == 45 & pix_y == 269)| (pix_x == 45 & pix_y == 270)| (pix_x == 45 & pix_y == 271)| (pix_x == 45 & pix_y == 272)| (pix_x == 45 & pix_y == 273)| (pix_x == 45 & pix_y == 294)| (pix_x == 45 & pix_y == 302)| (pix_x == 45 & pix_y == 303)| (pix_x == 45 & pix_y == 360)| (pix_x == 45 & pix_y == 361)| (pix_x == 45 & pix_y == 362)| (pix_x == 46 & pix_y == 252)| (pix_x == 46 & pix_y == 253)| (pix_x == 46 & pix_y == 266)| (pix_x == 46 & pix_y == 267)| (pix_x == 46 & pix_y == 268)| (pix_x == 46 & pix_y == 269)| (pix_x == 46 & pix_y == 270)| (pix_x == 46 & pix_y == 271)| (pix_x == 46 & pix_y == 294)| (pix_x == 47 & pix_y == 252)| (pix_x == 47 & pix_y == 253)| (pix_x == 47 & pix_y == 266)| (pix_x == 47 & pix_y == 267)| (pix_x == 47 & pix_y == 268)| (pix_x == 47 & pix_y == 269)| (pix_x == 47 & pix_y == 270)| (pix_x == 47 & pix_y == 271)| (pix_x == 47 & pix_y == 294)| (pix_x == 48 & pix_y == 351)| (pix_x == 48 & pix_y == 352)| (pix_x == 48 & pix_y == 363)| (pix_x == 48 & pix_y == 364)| (pix_x == 49 & pix_y == 351)| (pix_x == 49 & pix_y == 352)| (pix_x == 49 & pix_y == 363)| (pix_x == 49 & pix_y == 364)| (pix_x == 50 & pix_y == 363)| (pix_x == 50 & pix_y == 364)| (pix_x == 51 & pix_y == 363)| (pix_x == 51 & pix_y == 364)| (pix_x == 52 & pix_y == 363)| (pix_x == 52 & pix_y == 364)| (pix_x == 53 & pix_y == 341)| (pix_x == 53 & pix_y == 342)| (pix_x == 53 & pix_y == 343)| (pix_x == 53 & pix_y == 344)| (pix_x == 53 & pix_y == 345)| (pix_x == 53 & pix_y == 361)| (pix_x == 53 & pix_y == 362)| (pix_x == 53 & pix_y == 365)| (pix_x == 54 & pix_y == 341)| (pix_x == 54 & pix_y == 342)| (pix_x == 54 & pix_y == 343)| (pix_x == 54 & pix_y == 344)| (pix_x == 54 & pix_y == 345)| (pix_x == 54 & pix_y == 361)| (pix_x == 54 & pix_y == 362)| (pix_x == 54 & pix_y == 365)| (pix_x == 55 & pix_y == 360)| (pix_x == 55 & pix_y == 361)| (pix_x == 55 & pix_y == 362)| (pix_x == 55 & pix_y == 365)| (pix_x == 55 & pix_y == 369)| (pix_x == 55 & pix_y == 370)| (pix_x == 56 & pix_y == 360)| (pix_x == 56 & pix_y == 361)| (pix_x == 56 & pix_y == 362)| (pix_x == 56 & pix_y == 365)| (pix_x == 56 & pix_y == 369)| (pix_x == 56 & pix_y == 370)| (pix_x == 57 & pix_y == 360)| (pix_x == 57 & pix_y == 361)| (pix_x == 57 & pix_y == 362)| (pix_x == 57 & pix_y == 365)| (pix_x == 57 & pix_y == 369)| (pix_x == 57 & pix_y == 370)| (pix_x == 58 & pix_y == 353)| (pix_x == 58 & pix_y == 354)| (pix_x == 58 & pix_y == 361)| (pix_x == 58 & pix_y == 362)| (pix_x == 58 & pix_y == 363)| (pix_x == 58 & pix_y == 364)| (pix_x == 58 & pix_y == 368)| (pix_x == 59 & pix_y == 353)| (pix_x == 59 & pix_y == 354)| (pix_x == 59 & pix_y == 361)| (pix_x == 59 & pix_y == 362)| (pix_x == 59 & pix_y == 363)| (pix_x == 59 & pix_y == 364)| (pix_x == 59 & pix_y == 368)| (pix_x == 60 & pix_y == 345)| (pix_x == 60 & pix_y == 361)| (pix_x == 60 & pix_y == 362)| (pix_x == 60 & pix_y == 363)| (pix_x == 60 & pix_y == 364)| (pix_x == 60 & pix_y == 368)| (pix_x == 60 & pix_y == 369)| (pix_x == 60 & pix_y == 370)| (pix_x == 61 & pix_y == 345)| (pix_x == 61 & pix_y == 361)| (pix_x == 61 & pix_y == 362)| (pix_x == 61 & pix_y == 363)| (pix_x == 61 & pix_y == 364)| (pix_x == 61 & pix_y == 368)| (pix_x == 61 & pix_y == 369)| (pix_x == 61 & pix_y == 370)| (pix_x == 62 & pix_y == 360)| (pix_x == 62 & pix_y == 369)| (pix_x == 62 & pix_y == 370)| (pix_x == 63 & pix_y == 360)| (pix_x == 63 & pix_y == 369)| (pix_x == 63 & pix_y == 370)| (pix_x == 64 & pix_y == 360)| (pix_x == 64 & pix_y == 369)| (pix_x == 64 & pix_y == 370)| (pix_x == 65 & pix_y == 284)| (pix_x == 65 & pix_y == 338)| (pix_x == 65 & pix_y == 339)| (pix_x == 65 & pix_y == 356)| (pix_x == 65 & pix_y == 357)| (pix_x == 65 & pix_y == 358)| (pix_x == 65 & pix_y == 359)| (pix_x == 65 & pix_y == 361)| (pix_x == 65 & pix_y == 362)| (pix_x == 65 & pix_y == 366)| (pix_x == 65 & pix_y == 367)| (pix_x == 65 & pix_y == 368)| (pix_x == 65 & pix_y == 369)| (pix_x == 65 & pix_y == 370)| (pix_x == 65 & pix_y == 376)| (pix_x == 65 & pix_y == 377)| (pix_x == 66 & pix_y == 284)| (pix_x == 66 & pix_y == 338)| (pix_x == 66 & pix_y == 339)| (pix_x == 66 & pix_y == 356)| (pix_x == 66 & pix_y == 357)| (pix_x == 66 & pix_y == 358)| (pix_x == 66 & pix_y == 359)| (pix_x == 66 & pix_y == 361)| (pix_x == 66 & pix_y == 362)| (pix_x == 66 & pix_y == 366)| (pix_x == 66 & pix_y == 367)| (pix_x == 66 & pix_y == 368)| (pix_x == 66 & pix_y == 369)| (pix_x == 66 & pix_y == 370)| (pix_x == 66 & pix_y == 376)| (pix_x == 66 & pix_y == 377)| (pix_x == 67 & pix_y == 336)| (pix_x == 67 & pix_y == 337)| (pix_x == 67 & pix_y == 356)| (pix_x == 67 & pix_y == 357)| (pix_x == 67 & pix_y == 371)| (pix_x == 67 & pix_y == 372)| (pix_x == 68 & pix_y == 336)| (pix_x == 68 & pix_y == 337)| (pix_x == 68 & pix_y == 356)| (pix_x == 68 & pix_y == 357)| (pix_x == 68 & pix_y == 371)| (pix_x == 68 & pix_y == 372)| (pix_x == 69 & pix_y == 336)| (pix_x == 69 & pix_y == 337)| (pix_x == 69 & pix_y == 356)| (pix_x == 69 & pix_y == 357)| (pix_x == 69 & pix_y == 371)| (pix_x == 69 & pix_y == 372)| (pix_x == 70 & pix_y == 341)| (pix_x == 70 & pix_y == 342)| (pix_x == 70 & pix_y == 343)| (pix_x == 70 & pix_y == 344)| (pix_x == 70 & pix_y == 371)| (pix_x == 70 & pix_y == 372)| (pix_x == 71 & pix_y == 341)| (pix_x == 71 & pix_y == 342)| (pix_x == 71 & pix_y == 343)| (pix_x == 71 & pix_y == 344)| (pix_x == 71 & pix_y == 371)| (pix_x == 71 & pix_y == 372)| (pix_x == 72 & pix_y == 259)| (pix_x == 72 & pix_y == 260)| (pix_x == 72 & pix_y == 261)| (pix_x == 72 & pix_y == 343)| (pix_x == 72 & pix_y == 344)| (pix_x == 72 & pix_y == 345)| (pix_x == 72 & pix_y == 346)| (pix_x == 72 & pix_y == 347)| (pix_x == 72 & pix_y == 348)| (pix_x == 72 & pix_y == 349)| (pix_x == 72 & pix_y == 350)| (pix_x == 72 & pix_y == 361)| (pix_x == 72 & pix_y == 362)| (pix_x == 72 & pix_y == 371)| (pix_x == 72 & pix_y == 372)| (pix_x == 73 & pix_y == 259)| (pix_x == 73 & pix_y == 260)| (pix_x == 73 & pix_y == 261)| (pix_x == 73 & pix_y == 343)| (pix_x == 73 & pix_y == 344)| (pix_x == 73 & pix_y == 345)| (pix_x == 73 & pix_y == 346)| (pix_x == 73 & pix_y == 347)| (pix_x == 73 & pix_y == 348)| (pix_x == 73 & pix_y == 349)| (pix_x == 73 & pix_y == 350)| (pix_x == 73 & pix_y == 361)| (pix_x == 73 & pix_y == 362)| (pix_x == 73 & pix_y == 371)| (pix_x == 73 & pix_y == 372)| (pix_x == 74 & pix_y == 345)| (pix_x == 74 & pix_y == 346)| (pix_x == 74 & pix_y == 347)| (pix_x == 74 & pix_y == 348)| (pix_x == 74 & pix_y == 349)| (pix_x == 74 & pix_y == 361)| (pix_x == 74 & pix_y == 362)| (pix_x == 75 & pix_y == 345)| (pix_x == 75 & pix_y == 346)| (pix_x == 75 & pix_y == 347)| (pix_x == 75 & pix_y == 348)| (pix_x == 75 & pix_y == 349)| (pix_x == 75 & pix_y == 361)| (pix_x == 75 & pix_y == 362)| (pix_x == 76 & pix_y == 345)| (pix_x == 76 & pix_y == 346)| (pix_x == 76 & pix_y == 347)| (pix_x == 76 & pix_y == 348)| (pix_x == 76 & pix_y == 349)| (pix_x == 76 & pix_y == 361)| (pix_x == 76 & pix_y == 362)| (pix_x == 77 & pix_y == 351)| (pix_x == 77 & pix_y == 352)| (pix_x == 77 & pix_y == 373)| (pix_x == 77 & pix_y == 374)| (pix_x == 77 & pix_y == 375)| (pix_x == 78 & pix_y == 351)| (pix_x == 78 & pix_y == 352)| (pix_x == 78 & pix_y == 373)| (pix_x == 78 & pix_y == 374)| (pix_x == 78 & pix_y == 375)| (pix_x == 79 & pix_y == 251)| (pix_x == 79 & pix_y == 318)| (pix_x == 79 & pix_y == 319)| (pix_x == 79 & pix_y == 371)| (pix_x == 79 & pix_y == 372)| (pix_x == 79 & pix_y == 386)| (pix_x == 79 & pix_y == 387)| (pix_x == 79 & pix_y == 388)| (pix_x == 79 & pix_y == 389)| (pix_x == 79 & pix_y == 390)| (pix_x == 80 & pix_y == 251)| (pix_x == 80 & pix_y == 318)| (pix_x == 80 & pix_y == 319)| (pix_x == 80 & pix_y == 371)| (pix_x == 80 & pix_y == 372)| (pix_x == 80 & pix_y == 386)| (pix_x == 80 & pix_y == 387)| (pix_x == 80 & pix_y == 388)| (pix_x == 80 & pix_y == 389)| (pix_x == 80 & pix_y == 390)| (pix_x == 81 & pix_y == 251)| (pix_x == 81 & pix_y == 318)| (pix_x == 81 & pix_y == 319)| (pix_x == 81 & pix_y == 371)| (pix_x == 81 & pix_y == 372)| (pix_x == 81 & pix_y == 386)| (pix_x == 81 & pix_y == 387)| (pix_x == 81 & pix_y == 388)| (pix_x == 81 & pix_y == 389)| (pix_x == 81 & pix_y == 390)| (pix_x == 82 & pix_y == 310)| (pix_x == 82 & pix_y == 311)| (pix_x == 82 & pix_y == 355)| (pix_x == 82 & pix_y == 369)| (pix_x == 82 & pix_y == 370)| (pix_x == 82 & pix_y == 371)| (pix_x == 82 & pix_y == 372)| (pix_x == 82 & pix_y == 386)| (pix_x == 82 & pix_y == 387)| (pix_x == 82 & pix_y == 389)| (pix_x == 82 & pix_y == 390)| (pix_x == 83 & pix_y == 310)| (pix_x == 83 & pix_y == 311)| (pix_x == 83 & pix_y == 355)| (pix_x == 83 & pix_y == 369)| (pix_x == 83 & pix_y == 370)| (pix_x == 83 & pix_y == 371)| (pix_x == 83 & pix_y == 372)| (pix_x == 83 & pix_y == 386)| (pix_x == 83 & pix_y == 387)| (pix_x == 83 & pix_y == 389)| (pix_x == 83 & pix_y == 390)| (pix_x == 84 & pix_y == 282)| (pix_x == 84 & pix_y == 283)| (pix_x == 85 & pix_y == 282)| (pix_x == 85 & pix_y == 283)| (pix_x == 86 & pix_y == 313)| (pix_x == 86 & pix_y == 314)| (pix_x == 86 & pix_y == 406)| (pix_x == 87 & pix_y == 313)| (pix_x == 87 & pix_y == 314)| (pix_x == 87 & pix_y == 406)| (pix_x == 88 & pix_y == 313)| (pix_x == 88 & pix_y == 314)| (pix_x == 88 & pix_y == 406)| (pix_x == 89 & pix_y == 231)| (pix_x == 89 & pix_y == 232)| (pix_x == 89 & pix_y == 252)| (pix_x == 89 & pix_y == 253)| (pix_x == 89 & pix_y == 254)| (pix_x == 89 & pix_y == 255)| (pix_x == 89 & pix_y == 305)| (pix_x == 89 & pix_y == 306)| (pix_x == 89 & pix_y == 308)| (pix_x == 89 & pix_y == 309)| (pix_x == 89 & pix_y == 318)| (pix_x == 89 & pix_y == 319)| (pix_x == 90 & pix_y == 231)| (pix_x == 90 & pix_y == 232)| (pix_x == 90 & pix_y == 252)| (pix_x == 90 & pix_y == 253)| (pix_x == 90 & pix_y == 254)| (pix_x == 90 & pix_y == 255)| (pix_x == 90 & pix_y == 305)| (pix_x == 90 & pix_y == 306)| (pix_x == 90 & pix_y == 308)| (pix_x == 90 & pix_y == 309)| (pix_x == 90 & pix_y == 318)| (pix_x == 90 & pix_y == 319)| (pix_x == 91 & pix_y == 231)| (pix_x == 91 & pix_y == 232)| (pix_x == 91 & pix_y == 233)| (pix_x == 91 & pix_y == 292)| (pix_x == 91 & pix_y == 293)| (pix_x == 91 & pix_y == 318)| (pix_x == 91 & pix_y == 319)| (pix_x == 92 & pix_y == 231)| (pix_x == 92 & pix_y == 232)| (pix_x == 92 & pix_y == 233)| (pix_x == 92 & pix_y == 292)| (pix_x == 92 & pix_y == 293)| (pix_x == 92 & pix_y == 318)| (pix_x == 92 & pix_y == 319)| (pix_x == 93 & pix_y == 231)| (pix_x == 93 & pix_y == 232)| (pix_x == 93 & pix_y == 233)| (pix_x == 93 & pix_y == 292)| (pix_x == 93 & pix_y == 293)| (pix_x == 93 & pix_y == 318)| (pix_x == 93 & pix_y == 319)| (pix_x == 94 & pix_y == 402)| (pix_x == 94 & pix_y == 403)| (pix_x == 94 & pix_y == 409)| (pix_x == 94 & pix_y == 410)| (pix_x == 94 & pix_y == 412)| (pix_x == 94 & pix_y == 413)| (pix_x == 95 & pix_y == 402)| (pix_x == 95 & pix_y == 403)| (pix_x == 95 & pix_y == 409)| (pix_x == 95 & pix_y == 410)| (pix_x == 95 & pix_y == 412)| (pix_x == 95 & pix_y == 413)| (pix_x == 96 & pix_y == 239)| (pix_x == 96 & pix_y == 240)| (pix_x == 96 & pix_y == 241)| (pix_x == 96 & pix_y == 282)| (pix_x == 96 & pix_y == 283)| (pix_x == 96 & pix_y == 346)| (pix_x == 96 & pix_y == 347)| (pix_x == 96 & pix_y == 350)| (pix_x == 96 & pix_y == 371)| (pix_x == 96 & pix_y == 372)| (pix_x == 96 & pix_y == 384)| (pix_x == 96 & pix_y == 385)| (pix_x == 96 & pix_y == 412)| (pix_x == 96 & pix_y == 413)| (pix_x == 96 & pix_y == 431)| (pix_x == 97 & pix_y == 239)| (pix_x == 97 & pix_y == 240)| (pix_x == 97 & pix_y == 241)| (pix_x == 97 & pix_y == 282)| (pix_x == 97 & pix_y == 283)| (pix_x == 97 & pix_y == 346)| (pix_x == 97 & pix_y == 347)| (pix_x == 97 & pix_y == 350)| (pix_x == 97 & pix_y == 371)| (pix_x == 97 & pix_y == 372)| (pix_x == 97 & pix_y == 384)| (pix_x == 97 & pix_y == 385)| (pix_x == 97 & pix_y == 412)| (pix_x == 97 & pix_y == 413)| (pix_x == 97 & pix_y == 431)| (pix_x == 98 & pix_y == 224)| (pix_x == 98 & pix_y == 225)| (pix_x == 98 & pix_y == 310)| (pix_x == 98 & pix_y == 311)| (pix_x == 98 & pix_y == 312)| (pix_x == 98 & pix_y == 313)| (pix_x == 98 & pix_y == 314)| (pix_x == 98 & pix_y == 368)| (pix_x == 98 & pix_y == 419)| (pix_x == 98 & pix_y == 420)| (pix_x == 98 & pix_y == 421)| (pix_x == 99 & pix_y == 224)| (pix_x == 99 & pix_y == 225)| (pix_x == 99 & pix_y == 310)| (pix_x == 99 & pix_y == 311)| (pix_x == 99 & pix_y == 312)| (pix_x == 99 & pix_y == 313)| (pix_x == 99 & pix_y == 314)| (pix_x == 99 & pix_y == 368)| (pix_x == 99 & pix_y == 419)| (pix_x == 99 & pix_y == 420)| (pix_x == 99 & pix_y == 421)| (pix_x == 100 & pix_y == 224)| (pix_x == 100 & pix_y == 225)| (pix_x == 100 & pix_y == 310)| (pix_x == 100 & pix_y == 311)| (pix_x == 100 & pix_y == 312)| (pix_x == 100 & pix_y == 313)| (pix_x == 100 & pix_y == 314)| (pix_x == 100 & pix_y == 368)| (pix_x == 100 & pix_y == 419)| (pix_x == 100 & pix_y == 420)| (pix_x == 100 & pix_y == 421)| (pix_x == 101 & pix_y == 224)| (pix_x == 101 & pix_y == 225)| (pix_x == 101 & pix_y == 282)| (pix_x == 101 & pix_y == 283)| (pix_x == 101 & pix_y == 313)| (pix_x == 101 & pix_y == 314)| (pix_x == 101 & pix_y == 356)| (pix_x == 101 & pix_y == 357)| (pix_x == 101 & pix_y == 391)| (pix_x == 101 & pix_y == 392)| (pix_x == 101 & pix_y == 434)| (pix_x == 102 & pix_y == 224)| (pix_x == 102 & pix_y == 225)| (pix_x == 102 & pix_y == 282)| (pix_x == 102 & pix_y == 283)| (pix_x == 102 & pix_y == 313)| (pix_x == 102 & pix_y == 314)| (pix_x == 102 & pix_y == 356)| (pix_x == 102 & pix_y == 357)| (pix_x == 102 & pix_y == 391)| (pix_x == 102 & pix_y == 392)| (pix_x == 102 & pix_y == 434)| (pix_x == 103 & pix_y == 287)| (pix_x == 103 & pix_y == 288)| (pix_x == 103 & pix_y == 313)| (pix_x == 103 & pix_y == 314)| (pix_x == 103 & pix_y == 374)| (pix_x == 103 & pix_y == 375)| (pix_x == 103 & pix_y == 434)| (pix_x == 104 & pix_y == 287)| (pix_x == 104 & pix_y == 288)| (pix_x == 104 & pix_y == 313)| (pix_x == 104 & pix_y == 314)| (pix_x == 104 & pix_y == 374)| (pix_x == 104 & pix_y == 375)| (pix_x == 104 & pix_y == 434)| (pix_x == 105 & pix_y == 287)| (pix_x == 105 & pix_y == 288)| (pix_x == 105 & pix_y == 313)| (pix_x == 105 & pix_y == 314)| (pix_x == 105 & pix_y == 374)| (pix_x == 105 & pix_y == 375)| (pix_x == 105 & pix_y == 434)| (pix_x == 106 & pix_y == 355)| (pix_x == 107 & pix_y == 355)| (pix_x == 108 & pix_y == 261)| (pix_x == 108 & pix_y == 351)| (pix_x == 108 & pix_y == 352)| (pix_x == 109 & pix_y == 261)| (pix_x == 109 & pix_y == 351)| (pix_x == 109 & pix_y == 352)| (pix_x == 110 & pix_y == 277)| (pix_x == 110 & pix_y == 278)| (pix_x == 110 & pix_y == 279)| (pix_x == 110 & pix_y == 381)| (pix_x == 110 & pix_y == 382)| (pix_x == 111 & pix_y == 277)| (pix_x == 111 & pix_y == 278)| (pix_x == 111 & pix_y == 279)| (pix_x == 111 & pix_y == 381)| (pix_x == 111 & pix_y == 382)| (pix_x == 112 & pix_y == 277)| (pix_x == 112 & pix_y == 278)| (pix_x == 112 & pix_y == 279)| (pix_x == 112 & pix_y == 381)| (pix_x == 112 & pix_y == 382)| (pix_x == 113 & pix_y == 267)| (pix_x == 113 & pix_y == 268)| (pix_x == 113 & pix_y == 282)| (pix_x == 113 & pix_y == 283)| (pix_x == 113 & pix_y == 346)| (pix_x == 113 & pix_y == 347)| (pix_x == 114 & pix_y == 267)| (pix_x == 114 & pix_y == 268)| (pix_x == 114 & pix_y == 282)| (pix_x == 114 & pix_y == 283)| (pix_x == 114 & pix_y == 346)| (pix_x == 114 & pix_y == 347)| (pix_x == 115 & pix_y == 216)| (pix_x == 115 & pix_y == 217)| (pix_x == 115 & pix_y == 360)| (pix_x == 116 & pix_y == 216)| (pix_x == 116 & pix_y == 217)| (pix_x == 116 & pix_y == 360)| (pix_x == 117 & pix_y == 216)| (pix_x == 117 & pix_y == 217)| (pix_x == 117 & pix_y == 360)| (pix_x == 118 & pix_y == 351)| (pix_x == 118 & pix_y == 352)| (pix_x == 119 & pix_y == 351)| (pix_x == 119 & pix_y == 352)| (pix_x == 120 & pix_y == 315)| (pix_x == 120 & pix_y == 316)| (pix_x == 120 & pix_y == 356)| (pix_x == 120 & pix_y == 357)| (pix_x == 120 & pix_y == 358)| (pix_x == 120 & pix_y == 359)| (pix_x == 120 & pix_y == 417)| (pix_x == 120 & pix_y == 418)| (pix_x == 121 & pix_y == 315)| (pix_x == 121 & pix_y == 316)| (pix_x == 121 & pix_y == 356)| (pix_x == 121 & pix_y == 357)| (pix_x == 121 & pix_y == 358)| (pix_x == 121 & pix_y == 359)| (pix_x == 121 & pix_y == 417)| (pix_x == 121 & pix_y == 418)| (pix_x == 125 & pix_y == 211)| (pix_x == 125 & pix_y == 212)| (pix_x == 125 & pix_y == 219)| (pix_x == 125 & pix_y == 220)| (pix_x == 125 & pix_y == 221)| (pix_x == 125 & pix_y == 222)| (pix_x == 125 & pix_y == 238)| (pix_x == 125 & pix_y == 310)| (pix_x == 125 & pix_y == 311)| (pix_x == 125 & pix_y == 333)| (pix_x == 125 & pix_y == 334)| (pix_x == 126 & pix_y == 211)| (pix_x == 126 & pix_y == 212)| (pix_x == 126 & pix_y == 219)| (pix_x == 126 & pix_y == 220)| (pix_x == 126 & pix_y == 221)| (pix_x == 126 & pix_y == 222)| (pix_x == 126 & pix_y == 238)| (pix_x == 126 & pix_y == 310)| (pix_x == 126 & pix_y == 311)| (pix_x == 126 & pix_y == 333)| (pix_x == 126 & pix_y == 334)| (pix_x == 127 & pix_y == 228)| (pix_x == 127 & pix_y == 305)| (pix_x == 127 & pix_y == 306)| (pix_x == 127 & pix_y == 317)| (pix_x == 127 & pix_y == 318)| (pix_x == 127 & pix_y == 319)| (pix_x == 127 & pix_y == 335)| (pix_x == 128 & pix_y == 228)| (pix_x == 128 & pix_y == 305)| (pix_x == 128 & pix_y == 306)| (pix_x == 128 & pix_y == 317)| (pix_x == 128 & pix_y == 318)| (pix_x == 128 & pix_y == 319)| (pix_x == 128 & pix_y == 335)| (pix_x == 129 & pix_y == 228)| (pix_x == 129 & pix_y == 305)| (pix_x == 129 & pix_y == 306)| (pix_x == 129 & pix_y == 317)| (pix_x == 129 & pix_y == 318)| (pix_x == 129 & pix_y == 319)| (pix_x == 129 & pix_y == 335)| (pix_x == 130 & pix_y == 318)| (pix_x == 130 & pix_y == 319)| (pix_x == 130 & pix_y == 323)| (pix_x == 130 & pix_y == 324)| (pix_x == 130 & pix_y == 333)| (pix_x == 130 & pix_y == 334)| (pix_x == 130 & pix_y == 422)| (pix_x == 130 & pix_y == 423)| (pix_x == 130 & pix_y == 424)| (pix_x == 130 & pix_y == 425)| (pix_x == 131 & pix_y == 318)| (pix_x == 131 & pix_y == 319)| (pix_x == 131 & pix_y == 323)| (pix_x == 131 & pix_y == 324)| (pix_x == 131 & pix_y == 333)| (pix_x == 131 & pix_y == 334)| (pix_x == 131 & pix_y == 422)| (pix_x == 131 & pix_y == 423)| (pix_x == 131 & pix_y == 424)| (pix_x == 131 & pix_y == 425)| (pix_x == 132 & pix_y == 241)| (pix_x == 132 & pix_y == 257)| (pix_x == 132 & pix_y == 258)| (pix_x == 132 & pix_y == 264)| (pix_x == 132 & pix_y == 265)| (pix_x == 132 & pix_y == 312)| (pix_x == 132 & pix_y == 313)| (pix_x == 132 & pix_y == 314)| (pix_x == 132 & pix_y == 315)| (pix_x == 132 & pix_y == 316)| (pix_x == 132 & pix_y == 317)| (pix_x == 132 & pix_y == 318)| (pix_x == 132 & pix_y == 319)| (pix_x == 132 & pix_y == 345)| (pix_x == 133 & pix_y == 241)| (pix_x == 133 & pix_y == 257)| (pix_x == 133 & pix_y == 258)| (pix_x == 133 & pix_y == 264)| (pix_x == 133 & pix_y == 265)| (pix_x == 133 & pix_y == 312)| (pix_x == 133 & pix_y == 313)| (pix_x == 133 & pix_y == 314)| (pix_x == 133 & pix_y == 315)| (pix_x == 133 & pix_y == 316)| (pix_x == 133 & pix_y == 317)| (pix_x == 133 & pix_y == 318)| (pix_x == 133 & pix_y == 319)| (pix_x == 133 & pix_y == 345)| (pix_x == 134 & pix_y == 295)| (pix_x == 134 & pix_y == 296)| (pix_x == 134 & pix_y == 300)| (pix_x == 134 & pix_y == 301)| (pix_x == 134 & pix_y == 315)| (pix_x == 134 & pix_y == 316)| (pix_x == 134 & pix_y == 343)| (pix_x == 134 & pix_y == 344)| (pix_x == 134 & pix_y == 345)| (pix_x == 134 & pix_y == 346)| (pix_x == 134 & pix_y == 347)| (pix_x == 134 & pix_y == 426)| (pix_x == 135 & pix_y == 295)| (pix_x == 135 & pix_y == 296)| (pix_x == 135 & pix_y == 300)| (pix_x == 135 & pix_y == 301)| (pix_x == 135 & pix_y == 315)| (pix_x == 135 & pix_y == 316)| (pix_x == 135 & pix_y == 343)| (pix_x == 135 & pix_y == 344)| (pix_x == 135 & pix_y == 345)| (pix_x == 135 & pix_y == 346)| (pix_x == 135 & pix_y == 347)| (pix_x == 135 & pix_y == 426)| (pix_x == 136 & pix_y == 295)| (pix_x == 136 & pix_y == 296)| (pix_x == 136 & pix_y == 300)| (pix_x == 136 & pix_y == 301)| (pix_x == 136 & pix_y == 315)| (pix_x == 136 & pix_y == 316)| (pix_x == 136 & pix_y == 343)| (pix_x == 136 & pix_y == 344)| (pix_x == 136 & pix_y == 345)| (pix_x == 136 & pix_y == 346)| (pix_x == 136 & pix_y == 347)| (pix_x == 136 & pix_y == 426)| (pix_x == 137 & pix_y == 206)| (pix_x == 137 & pix_y == 207)| (pix_x == 137 & pix_y == 209)| (pix_x == 137 & pix_y == 210)| (pix_x == 137 & pix_y == 262)| (pix_x == 137 & pix_y == 263)| (pix_x == 137 & pix_y == 264)| (pix_x == 137 & pix_y == 265)| (pix_x == 137 & pix_y == 302)| (pix_x == 137 & pix_y == 303)| (pix_x == 137 & pix_y == 304)| (pix_x == 137 & pix_y == 310)| (pix_x == 137 & pix_y == 311)| (pix_x == 137 & pix_y == 312)| (pix_x == 137 & pix_y == 313)| (pix_x == 137 & pix_y == 314)| (pix_x == 137 & pix_y == 345)| (pix_x == 137 & pix_y == 346)| (pix_x == 137 & pix_y == 347)| (pix_x == 137 & pix_y == 426)| (pix_x == 138 & pix_y == 206)| (pix_x == 138 & pix_y == 207)| (pix_x == 138 & pix_y == 209)| (pix_x == 138 & pix_y == 210)| (pix_x == 138 & pix_y == 262)| (pix_x == 138 & pix_y == 263)| (pix_x == 138 & pix_y == 264)| (pix_x == 138 & pix_y == 265)| (pix_x == 138 & pix_y == 302)| (pix_x == 138 & pix_y == 303)| (pix_x == 138 & pix_y == 304)| (pix_x == 138 & pix_y == 310)| (pix_x == 138 & pix_y == 311)| (pix_x == 138 & pix_y == 312)| (pix_x == 138 & pix_y == 313)| (pix_x == 138 & pix_y == 314)| (pix_x == 138 & pix_y == 345)| (pix_x == 138 & pix_y == 346)| (pix_x == 138 & pix_y == 347)| (pix_x == 138 & pix_y == 426)| (pix_x == 139 & pix_y == 206)| (pix_x == 139 & pix_y == 207)| (pix_x == 139 & pix_y == 257)| (pix_x == 139 & pix_y == 258)| (pix_x == 139 & pix_y == 264)| (pix_x == 139 & pix_y == 265)| (pix_x == 139 & pix_y == 343)| (pix_x == 139 & pix_y == 344)| (pix_x == 139 & pix_y == 345)| (pix_x == 139 & pix_y == 346)| (pix_x == 139 & pix_y == 347)| (pix_x == 139 & pix_y == 350)| (pix_x == 139 & pix_y == 351)| (pix_x == 139 & pix_y == 352)| (pix_x == 140 & pix_y == 206)| (pix_x == 140 & pix_y == 207)| (pix_x == 140 & pix_y == 257)| (pix_x == 140 & pix_y == 258)| (pix_x == 140 & pix_y == 264)| (pix_x == 140 & pix_y == 265)| (pix_x == 140 & pix_y == 343)| (pix_x == 140 & pix_y == 344)| (pix_x == 140 & pix_y == 345)| (pix_x == 140 & pix_y == 346)| (pix_x == 140 & pix_y == 347)| (pix_x == 140 & pix_y == 350)| (pix_x == 140 & pix_y == 351)| (pix_x == 140 & pix_y == 352)| (pix_x == 141 & pix_y == 206)| (pix_x == 141 & pix_y == 207)| (pix_x == 141 & pix_y == 257)| (pix_x == 141 & pix_y == 258)| (pix_x == 141 & pix_y == 264)| (pix_x == 141 & pix_y == 265)| (pix_x == 141 & pix_y == 343)| (pix_x == 141 & pix_y == 344)| (pix_x == 141 & pix_y == 345)| (pix_x == 141 & pix_y == 346)| (pix_x == 141 & pix_y == 347)| (pix_x == 141 & pix_y == 350)| (pix_x == 141 & pix_y == 351)| (pix_x == 141 & pix_y == 352)| (pix_x == 142 & pix_y == 198)| (pix_x == 142 & pix_y == 199)| (pix_x == 142 & pix_y == 200)| (pix_x == 142 & pix_y == 228)| (pix_x == 142 & pix_y == 264)| (pix_x == 142 & pix_y == 265)| (pix_x == 142 & pix_y == 266)| (pix_x == 142 & pix_y == 302)| (pix_x == 142 & pix_y == 303)| (pix_x == 142 & pix_y == 312)| (pix_x == 142 & pix_y == 313)| (pix_x == 142 & pix_y == 314)| (pix_x == 142 & pix_y == 323)| (pix_x == 142 & pix_y == 324)| (pix_x == 142 & pix_y == 348)| (pix_x == 142 & pix_y == 349)| (pix_x == 143 & pix_y == 198)| (pix_x == 143 & pix_y == 199)| (pix_x == 143 & pix_y == 200)| (pix_x == 143 & pix_y == 228)| (pix_x == 143 & pix_y == 264)| (pix_x == 143 & pix_y == 265)| (pix_x == 143 & pix_y == 266)| (pix_x == 143 & pix_y == 302)| (pix_x == 143 & pix_y == 303)| (pix_x == 143 & pix_y == 312)| (pix_x == 143 & pix_y == 313)| (pix_x == 143 & pix_y == 314)| (pix_x == 143 & pix_y == 323)| (pix_x == 143 & pix_y == 324)| (pix_x == 143 & pix_y == 348)| (pix_x == 143 & pix_y == 349)| (pix_x == 144 & pix_y == 251)| (pix_x == 144 & pix_y == 264)| (pix_x == 144 & pix_y == 265)| (pix_x == 144 & pix_y == 266)| (pix_x == 144 & pix_y == 302)| (pix_x == 144 & pix_y == 303)| (pix_x == 144 & pix_y == 348)| (pix_x == 144 & pix_y == 349)| (pix_x == 144 & pix_y == 350)| (pix_x == 144 & pix_y == 351)| (pix_x == 144 & pix_y == 352)| (pix_x == 144 & pix_y == 381)| (pix_x == 144 & pix_y == 382)| (pix_x == 144 & pix_y == 388)| (pix_x == 145 & pix_y == 251)| (pix_x == 145 & pix_y == 264)| (pix_x == 145 & pix_y == 265)| (pix_x == 145 & pix_y == 266)| (pix_x == 145 & pix_y == 302)| (pix_x == 145 & pix_y == 303)| (pix_x == 145 & pix_y == 348)| (pix_x == 145 & pix_y == 349)| (pix_x == 145 & pix_y == 350)| (pix_x == 145 & pix_y == 351)| (pix_x == 145 & pix_y == 352)| (pix_x == 145 & pix_y == 381)| (pix_x == 145 & pix_y == 382)| (pix_x == 145 & pix_y == 388)| (pix_x == 146 & pix_y == 262)| (pix_x == 146 & pix_y == 263)| (pix_x == 146 & pix_y == 264)| (pix_x == 146 & pix_y == 265)| (pix_x == 146 & pix_y == 289)| (pix_x == 146 & pix_y == 302)| (pix_x == 146 & pix_y == 303)| (pix_x == 146 & pix_y == 341)| (pix_x == 146 & pix_y == 342)| (pix_x == 146 & pix_y == 388)| (pix_x == 147 & pix_y == 262)| (pix_x == 147 & pix_y == 263)| (pix_x == 147 & pix_y == 264)| (pix_x == 147 & pix_y == 265)| (pix_x == 147 & pix_y == 289)| (pix_x == 147 & pix_y == 302)| (pix_x == 147 & pix_y == 303)| (pix_x == 147 & pix_y == 341)| (pix_x == 147 & pix_y == 342)| (pix_x == 147 & pix_y == 388)| (pix_x == 148 & pix_y == 262)| (pix_x == 148 & pix_y == 263)| (pix_x == 148 & pix_y == 264)| (pix_x == 148 & pix_y == 265)| (pix_x == 148 & pix_y == 289)| (pix_x == 148 & pix_y == 302)| (pix_x == 148 & pix_y == 303)| (pix_x == 148 & pix_y == 341)| (pix_x == 148 & pix_y == 342)| (pix_x == 148 & pix_y == 388)| (pix_x == 149 & pix_y == 241)| (pix_x == 149 & pix_y == 259)| (pix_x == 149 & pix_y == 260)| (pix_x == 149 & pix_y == 264)| (pix_x == 149 & pix_y == 265)| (pix_x == 149 & pix_y == 269)| (pix_x == 149 & pix_y == 270)| (pix_x == 149 & pix_y == 271)| (pix_x == 149 & pix_y == 277)| (pix_x == 149 & pix_y == 278)| (pix_x == 149 & pix_y == 300)| (pix_x == 149 & pix_y == 301)| (pix_x == 149 & pix_y == 302)| (pix_x == 149 & pix_y == 303)| (pix_x == 149 & pix_y == 340)| (pix_x == 149 & pix_y == 341)| (pix_x == 149 & pix_y == 342)| (pix_x == 149 & pix_y == 353)| (pix_x == 149 & pix_y == 354)| (pix_x == 149 & pix_y == 356)| (pix_x == 149 & pix_y == 357)| (pix_x == 149 & pix_y == 445)| (pix_x == 149 & pix_y == 446)| (pix_x == 150 & pix_y == 241)| (pix_x == 150 & pix_y == 259)| (pix_x == 150 & pix_y == 260)| (pix_x == 150 & pix_y == 264)| (pix_x == 150 & pix_y == 265)| (pix_x == 150 & pix_y == 269)| (pix_x == 150 & pix_y == 270)| (pix_x == 150 & pix_y == 271)| (pix_x == 150 & pix_y == 277)| (pix_x == 150 & pix_y == 278)| (pix_x == 150 & pix_y == 300)| (pix_x == 150 & pix_y == 301)| (pix_x == 150 & pix_y == 302)| (pix_x == 150 & pix_y == 303)| (pix_x == 150 & pix_y == 340)| (pix_x == 150 & pix_y == 341)| (pix_x == 150 & pix_y == 342)| (pix_x == 150 & pix_y == 353)| (pix_x == 150 & pix_y == 354)| (pix_x == 150 & pix_y == 356)| (pix_x == 150 & pix_y == 357)| (pix_x == 150 & pix_y == 445)| (pix_x == 150 & pix_y == 446)| (pix_x == 151 & pix_y == 238)| (pix_x == 151 & pix_y == 269)| (pix_x == 151 & pix_y == 270)| (pix_x == 151 & pix_y == 271)| (pix_x == 151 & pix_y == 272)| (pix_x == 151 & pix_y == 273)| (pix_x == 151 & pix_y == 277)| (pix_x == 151 & pix_y == 278)| (pix_x == 151 & pix_y == 374)| (pix_x == 151 & pix_y == 375)| (pix_x == 152 & pix_y == 238)| (pix_x == 152 & pix_y == 269)| (pix_x == 152 & pix_y == 270)| (pix_x == 152 & pix_y == 271)| (pix_x == 152 & pix_y == 272)| (pix_x == 152 & pix_y == 273)| (pix_x == 152 & pix_y == 277)| (pix_x == 152 & pix_y == 278)| (pix_x == 152 & pix_y == 374)| (pix_x == 152 & pix_y == 375)| (pix_x == 153 & pix_y == 238)| (pix_x == 153 & pix_y == 269)| (pix_x == 153 & pix_y == 270)| (pix_x == 153 & pix_y == 271)| (pix_x == 153 & pix_y == 272)| (pix_x == 153 & pix_y == 273)| (pix_x == 153 & pix_y == 277)| (pix_x == 153 & pix_y == 278)| (pix_x == 153 & pix_y == 374)| (pix_x == 153 & pix_y == 375)| (pix_x == 154 & pix_y == 201)| (pix_x == 154 & pix_y == 202)| (pix_x == 154 & pix_y == 264)| (pix_x == 154 & pix_y == 265)| (pix_x == 154 & pix_y == 272)| (pix_x == 154 & pix_y == 273)| (pix_x == 154 & pix_y == 328)| (pix_x == 154 & pix_y == 329)| (pix_x == 154 & pix_y == 332)| (pix_x == 154 & pix_y == 355)| (pix_x == 154 & pix_y == 360)| (pix_x == 155 & pix_y == 201)| (pix_x == 155 & pix_y == 202)| (pix_x == 155 & pix_y == 264)| (pix_x == 155 & pix_y == 265)| (pix_x == 155 & pix_y == 272)| (pix_x == 155 & pix_y == 273)| (pix_x == 155 & pix_y == 328)| (pix_x == 155 & pix_y == 329)| (pix_x == 155 & pix_y == 332)| (pix_x == 155 & pix_y == 355)| (pix_x == 155 & pix_y == 360)| (pix_x == 156 & pix_y == 358)| (pix_x == 156 & pix_y == 359)| (pix_x == 156 & pix_y == 442)| (pix_x == 156 & pix_y == 443)| (pix_x == 157 & pix_y == 358)| (pix_x == 157 & pix_y == 359)| (pix_x == 157 & pix_y == 442)| (pix_x == 157 & pix_y == 443)| (pix_x == 158 & pix_y == 267)| (pix_x == 158 & pix_y == 268)| (pix_x == 158 & pix_y == 325)| (pix_x == 158 & pix_y == 326)| (pix_x == 158 & pix_y == 394)| (pix_x == 158 & pix_y == 395)| (pix_x == 158 & pix_y == 419)| (pix_x == 158 & pix_y == 420)| (pix_x == 158 & pix_y == 442)| (pix_x == 158 & pix_y == 443)| (pix_x == 158 & pix_y == 444)| (pix_x == 159 & pix_y == 267)| (pix_x == 159 & pix_y == 268)| (pix_x == 159 & pix_y == 325)| (pix_x == 159 & pix_y == 326)| (pix_x == 159 & pix_y == 394)| (pix_x == 159 & pix_y == 395)| (pix_x == 159 & pix_y == 419)| (pix_x == 159 & pix_y == 420)| (pix_x == 159 & pix_y == 442)| (pix_x == 159 & pix_y == 443)| (pix_x == 159 & pix_y == 444)| (pix_x == 160 & pix_y == 267)| (pix_x == 160 & pix_y == 268)| (pix_x == 160 & pix_y == 325)| (pix_x == 160 & pix_y == 326)| (pix_x == 160 & pix_y == 394)| (pix_x == 160 & pix_y == 395)| (pix_x == 160 & pix_y == 419)| (pix_x == 160 & pix_y == 420)| (pix_x == 160 & pix_y == 442)| (pix_x == 160 & pix_y == 443)| (pix_x == 160 & pix_y == 444)| (pix_x == 161 & pix_y == 323)| (pix_x == 161 & pix_y == 324)| (pix_x == 161 & pix_y == 356)| (pix_x == 161 & pix_y == 357)| (pix_x == 161 & pix_y == 388)| (pix_x == 161 & pix_y == 442)| (pix_x == 161 & pix_y == 443)| (pix_x == 162 & pix_y == 323)| (pix_x == 162 & pix_y == 324)| (pix_x == 162 & pix_y == 356)| (pix_x == 162 & pix_y == 357)| (pix_x == 162 & pix_y == 388)| (pix_x == 162 & pix_y == 442)| (pix_x == 162 & pix_y == 443)| (pix_x == 163 & pix_y == 317)| (pix_x == 163 & pix_y == 356)| (pix_x == 163 & pix_y == 357)| (pix_x == 163 & pix_y == 360)| (pix_x == 163 & pix_y == 402)| (pix_x == 163 & pix_y == 403)| (pix_x == 163 & pix_y == 437)| (pix_x == 163 & pix_y == 438)| (pix_x == 164 & pix_y == 317)| (pix_x == 164 & pix_y == 356)| (pix_x == 164 & pix_y == 357)| (pix_x == 164 & pix_y == 360)| (pix_x == 164 & pix_y == 402)| (pix_x == 164 & pix_y == 403)| (pix_x == 164 & pix_y == 437)| (pix_x == 164 & pix_y == 438)| (pix_x == 165 & pix_y == 317)| (pix_x == 165 & pix_y == 356)| (pix_x == 165 & pix_y == 357)| (pix_x == 165 & pix_y == 360)| (pix_x == 165 & pix_y == 402)| (pix_x == 165 & pix_y == 403)| (pix_x == 165 & pix_y == 437)| (pix_x == 165 & pix_y == 438)| (pix_x == 168 & pix_y == 369)| (pix_x == 168 & pix_y == 370)| (pix_x == 168 & pix_y == 388)| (pix_x == 169 & pix_y == 369)| (pix_x == 169 & pix_y == 370)| (pix_x == 169 & pix_y == 388)| (pix_x == 170 & pix_y == 264)| (pix_x == 170 & pix_y == 265)| (pix_x == 170 & pix_y == 266)| (pix_x == 170 & pix_y == 406)| (pix_x == 170 & pix_y == 431)| (pix_x == 170 & pix_y == 432)| (pix_x == 170 & pix_y == 433)| (pix_x == 170 & pix_y == 435)| (pix_x == 170 & pix_y == 436)| (pix_x == 171 & pix_y == 264)| (pix_x == 171 & pix_y == 265)| (pix_x == 171 & pix_y == 266)| (pix_x == 171 & pix_y == 406)| (pix_x == 171 & pix_y == 431)| (pix_x == 171 & pix_y == 432)| (pix_x == 171 & pix_y == 433)| (pix_x == 171 & pix_y == 435)| (pix_x == 171 & pix_y == 436)| (pix_x == 172 & pix_y == 264)| (pix_x == 172 & pix_y == 265)| (pix_x == 172 & pix_y == 266)| (pix_x == 172 & pix_y == 406)| (pix_x == 172 & pix_y == 431)| (pix_x == 172 & pix_y == 432)| (pix_x == 172 & pix_y == 433)| (pix_x == 172 & pix_y == 435)| (pix_x == 172 & pix_y == 436)| (pix_x == 173 & pix_y == 266)| (pix_x == 173 & pix_y == 275)| (pix_x == 173 & pix_y == 276)| (pix_x == 173 & pix_y == 297)| (pix_x == 173 & pix_y == 298)| (pix_x == 173 & pix_y == 386)| (pix_x == 173 & pix_y == 387)| (pix_x == 173 & pix_y == 391)| (pix_x == 173 & pix_y == 392)| (pix_x == 173 & pix_y == 402)| (pix_x == 173 & pix_y == 403)| (pix_x == 173 & pix_y == 432)| (pix_x == 173 & pix_y == 433)| (pix_x == 173 & pix_y == 434)| (pix_x == 173 & pix_y == 435)| (pix_x == 173 & pix_y == 436)| (pix_x == 173 & pix_y == 437)| (pix_x == 173 & pix_y == 438)| (pix_x == 173 & pix_y == 439)| (pix_x == 174 & pix_y == 266)| (pix_x == 174 & pix_y == 275)| (pix_x == 174 & pix_y == 276)| (pix_x == 174 & pix_y == 297)| (pix_x == 174 & pix_y == 298)| (pix_x == 174 & pix_y == 386)| (pix_x == 174 & pix_y == 387)| (pix_x == 174 & pix_y == 391)| (pix_x == 174 & pix_y == 392)| (pix_x == 174 & pix_y == 402)| (pix_x == 174 & pix_y == 403)| (pix_x == 174 & pix_y == 432)| (pix_x == 174 & pix_y == 433)| (pix_x == 174 & pix_y == 434)| (pix_x == 174 & pix_y == 435)| (pix_x == 174 & pix_y == 436)| (pix_x == 174 & pix_y == 437)| (pix_x == 174 & pix_y == 438)| (pix_x == 174 & pix_y == 439)| (pix_x == 175 & pix_y == 224)| (pix_x == 175 & pix_y == 225)| (pix_x == 175 & pix_y == 226)| (pix_x == 175 & pix_y == 227)| (pix_x == 175 & pix_y == 234)| (pix_x == 175 & pix_y == 235)| (pix_x == 175 & pix_y == 266)| (pix_x == 175 & pix_y == 295)| (pix_x == 175 & pix_y == 296)| (pix_x == 175 & pix_y == 384)| (pix_x == 175 & pix_y == 385)| (pix_x == 175 & pix_y == 386)| (pix_x == 175 & pix_y == 387)| (pix_x == 175 & pix_y == 402)| (pix_x == 175 & pix_y == 403)| (pix_x == 175 & pix_y == 406)| (pix_x == 175 & pix_y == 407)| (pix_x == 175 & pix_y == 408)| (pix_x == 175 & pix_y == 409)| (pix_x == 175 & pix_y == 410)| (pix_x == 175 & pix_y == 426)| (pix_x == 175 & pix_y == 432)| (pix_x == 175 & pix_y == 433)| (pix_x == 175 & pix_y == 434)| (pix_x == 175 & pix_y == 435)| (pix_x == 175 & pix_y == 436)| (pix_x == 175 & pix_y == 437)| (pix_x == 175 & pix_y == 438)| (pix_x == 175 & pix_y == 439)| (pix_x == 175 & pix_y == 440)| (pix_x == 175 & pix_y == 441)| (pix_x == 176 & pix_y == 224)| (pix_x == 176 & pix_y == 225)| (pix_x == 176 & pix_y == 226)| (pix_x == 176 & pix_y == 227)| (pix_x == 176 & pix_y == 234)| (pix_x == 176 & pix_y == 235)| (pix_x == 176 & pix_y == 266)| (pix_x == 176 & pix_y == 295)| (pix_x == 176 & pix_y == 296)| (pix_x == 176 & pix_y == 384)| (pix_x == 176 & pix_y == 385)| (pix_x == 176 & pix_y == 386)| (pix_x == 176 & pix_y == 387)| (pix_x == 176 & pix_y == 402)| (pix_x == 176 & pix_y == 403)| (pix_x == 176 & pix_y == 406)| (pix_x == 176 & pix_y == 407)| (pix_x == 176 & pix_y == 408)| (pix_x == 176 & pix_y == 409)| (pix_x == 176 & pix_y == 410)| (pix_x == 176 & pix_y == 426)| (pix_x == 176 & pix_y == 432)| (pix_x == 176 & pix_y == 433)| (pix_x == 176 & pix_y == 434)| (pix_x == 176 & pix_y == 435)| (pix_x == 176 & pix_y == 436)| (pix_x == 176 & pix_y == 437)| (pix_x == 176 & pix_y == 438)| (pix_x == 176 & pix_y == 439)| (pix_x == 176 & pix_y == 440)| (pix_x == 176 & pix_y == 441)| (pix_x == 177 & pix_y == 224)| (pix_x == 177 & pix_y == 225)| (pix_x == 177 & pix_y == 226)| (pix_x == 177 & pix_y == 227)| (pix_x == 177 & pix_y == 234)| (pix_x == 177 & pix_y == 235)| (pix_x == 177 & pix_y == 266)| (pix_x == 177 & pix_y == 295)| (pix_x == 177 & pix_y == 296)| (pix_x == 177 & pix_y == 384)| (pix_x == 177 & pix_y == 385)| (pix_x == 177 & pix_y == 386)| (pix_x == 177 & pix_y == 387)| (pix_x == 177 & pix_y == 402)| (pix_x == 177 & pix_y == 403)| (pix_x == 177 & pix_y == 406)| (pix_x == 177 & pix_y == 407)| (pix_x == 177 & pix_y == 408)| (pix_x == 177 & pix_y == 409)| (pix_x == 177 & pix_y == 410)| (pix_x == 177 & pix_y == 426)| (pix_x == 177 & pix_y == 432)| (pix_x == 177 & pix_y == 433)| (pix_x == 177 & pix_y == 434)| (pix_x == 177 & pix_y == 435)| (pix_x == 177 & pix_y == 436)| (pix_x == 177 & pix_y == 437)| (pix_x == 177 & pix_y == 438)| (pix_x == 177 & pix_y == 439)| (pix_x == 177 & pix_y == 440)| (pix_x == 177 & pix_y == 441)| (pix_x == 178 & pix_y == 196)| (pix_x == 178 & pix_y == 197)| (pix_x == 178 & pix_y == 200)| (pix_x == 178 & pix_y == 257)| (pix_x == 178 & pix_y == 258)| (pix_x == 178 & pix_y == 264)| (pix_x == 178 & pix_y == 265)| (pix_x == 178 & pix_y == 297)| (pix_x == 178 & pix_y == 298)| (pix_x == 178 & pix_y == 384)| (pix_x == 178 & pix_y == 385)| (pix_x == 178 & pix_y == 401)| (pix_x == 178 & pix_y == 406)| (pix_x == 178 & pix_y == 407)| (pix_x == 178 & pix_y == 408)| (pix_x == 178 & pix_y == 424)| (pix_x == 178 & pix_y == 425)| (pix_x == 178 & pix_y == 432)| (pix_x == 178 & pix_y == 433)| (pix_x == 178 & pix_y == 434)| (pix_x == 178 & pix_y == 435)| (pix_x == 178 & pix_y == 436)| (pix_x == 178 & pix_y == 437)| (pix_x == 178 & pix_y == 438)| (pix_x == 178 & pix_y == 439)| (pix_x == 178 & pix_y == 440)| (pix_x == 178 & pix_y == 441)| (pix_x == 179 & pix_y == 196)| (pix_x == 179 & pix_y == 197)| (pix_x == 179 & pix_y == 200)| (pix_x == 179 & pix_y == 257)| (pix_x == 179 & pix_y == 258)| (pix_x == 179 & pix_y == 264)| (pix_x == 179 & pix_y == 265)| (pix_x == 179 & pix_y == 297)| (pix_x == 179 & pix_y == 298)| (pix_x == 179 & pix_y == 384)| (pix_x == 179 & pix_y == 385)| (pix_x == 179 & pix_y == 401)| (pix_x == 179 & pix_y == 406)| (pix_x == 179 & pix_y == 407)| (pix_x == 179 & pix_y == 408)| (pix_x == 179 & pix_y == 424)| (pix_x == 179 & pix_y == 425)| (pix_x == 179 & pix_y == 432)| (pix_x == 179 & pix_y == 433)| (pix_x == 179 & pix_y == 434)| (pix_x == 179 & pix_y == 435)| (pix_x == 179 & pix_y == 436)| (pix_x == 179 & pix_y == 437)| (pix_x == 179 & pix_y == 438)| (pix_x == 179 & pix_y == 439)| (pix_x == 179 & pix_y == 440)| (pix_x == 179 & pix_y == 441)| (pix_x == 180 & pix_y == 196)| (pix_x == 180 & pix_y == 197)| (pix_x == 180 & pix_y == 198)| (pix_x == 180 & pix_y == 199)| (pix_x == 180 & pix_y == 200)| (pix_x == 180 & pix_y == 224)| (pix_x == 180 & pix_y == 225)| (pix_x == 180 & pix_y == 383)| (pix_x == 180 & pix_y == 399)| (pix_x == 180 & pix_y == 400)| (pix_x == 180 & pix_y == 401)| (pix_x == 180 & pix_y == 406)| (pix_x == 180 & pix_y == 434)| (pix_x == 180 & pix_y == 435)| (pix_x == 180 & pix_y == 436)| (pix_x == 180 & pix_y == 437)| (pix_x == 180 & pix_y == 438)| (pix_x == 181 & pix_y == 196)| (pix_x == 181 & pix_y == 197)| (pix_x == 181 & pix_y == 198)| (pix_x == 181 & pix_y == 199)| (pix_x == 181 & pix_y == 200)| (pix_x == 181 & pix_y == 224)| (pix_x == 181 & pix_y == 225)| (pix_x == 181 & pix_y == 383)| (pix_x == 181 & pix_y == 399)| (pix_x == 181 & pix_y == 400)| (pix_x == 181 & pix_y == 401)| (pix_x == 181 & pix_y == 406)| (pix_x == 181 & pix_y == 434)| (pix_x == 181 & pix_y == 435)| (pix_x == 181 & pix_y == 436)| (pix_x == 181 & pix_y == 437)| (pix_x == 181 & pix_y == 438)| (pix_x == 182 & pix_y == 196)| (pix_x == 182 & pix_y == 197)| (pix_x == 182 & pix_y == 206)| (pix_x == 182 & pix_y == 207)| (pix_x == 182 & pix_y == 208)| (pix_x == 182 & pix_y == 218)| (pix_x == 182 & pix_y == 219)| (pix_x == 182 & pix_y == 220)| (pix_x == 182 & pix_y == 223)| (pix_x == 182 & pix_y == 247)| (pix_x == 182 & pix_y == 248)| (pix_x == 182 & pix_y == 249)| (pix_x == 182 & pix_y == 250)| (pix_x == 182 & pix_y == 383)| (pix_x == 182 & pix_y == 384)| (pix_x == 182 & pix_y == 385)| (pix_x == 182 & pix_y == 432)| (pix_x == 182 & pix_y == 433)| (pix_x == 182 & pix_y == 434)| (pix_x == 182 & pix_y == 435)| (pix_x == 182 & pix_y == 436)| (pix_x == 182 & pix_y == 437)| (pix_x == 182 & pix_y == 438)| (pix_x == 183 & pix_y == 196)| (pix_x == 183 & pix_y == 197)| (pix_x == 183 & pix_y == 206)| (pix_x == 183 & pix_y == 207)| (pix_x == 183 & pix_y == 208)| (pix_x == 183 & pix_y == 218)| (pix_x == 183 & pix_y == 219)| (pix_x == 183 & pix_y == 220)| (pix_x == 183 & pix_y == 223)| (pix_x == 183 & pix_y == 247)| (pix_x == 183 & pix_y == 248)| (pix_x == 183 & pix_y == 249)| (pix_x == 183 & pix_y == 250)| (pix_x == 183 & pix_y == 383)| (pix_x == 183 & pix_y == 384)| (pix_x == 183 & pix_y == 385)| (pix_x == 183 & pix_y == 432)| (pix_x == 183 & pix_y == 433)| (pix_x == 183 & pix_y == 434)| (pix_x == 183 & pix_y == 435)| (pix_x == 183 & pix_y == 436)| (pix_x == 183 & pix_y == 437)| (pix_x == 183 & pix_y == 438)| (pix_x == 184 & pix_y == 196)| (pix_x == 184 & pix_y == 197)| (pix_x == 184 & pix_y == 206)| (pix_x == 184 & pix_y == 207)| (pix_x == 184 & pix_y == 208)| (pix_x == 184 & pix_y == 218)| (pix_x == 184 & pix_y == 219)| (pix_x == 184 & pix_y == 220)| (pix_x == 184 & pix_y == 223)| (pix_x == 184 & pix_y == 247)| (pix_x == 184 & pix_y == 248)| (pix_x == 184 & pix_y == 249)| (pix_x == 184 & pix_y == 250)| (pix_x == 184 & pix_y == 383)| (pix_x == 184 & pix_y == 384)| (pix_x == 184 & pix_y == 385)| (pix_x == 184 & pix_y == 432)| (pix_x == 184 & pix_y == 433)| (pix_x == 184 & pix_y == 434)| (pix_x == 184 & pix_y == 435)| (pix_x == 184 & pix_y == 436)| (pix_x == 184 & pix_y == 437)| (pix_x == 184 & pix_y == 438)| (pix_x == 185 & pix_y == 206)| (pix_x == 185 & pix_y == 207)| (pix_x == 185 & pix_y == 208)| (pix_x == 185 & pix_y == 251)| (pix_x == 185 & pix_y == 384)| (pix_x == 185 & pix_y == 385)| (pix_x == 185 & pix_y == 432)| (pix_x == 185 & pix_y == 433)| (pix_x == 185 & pix_y == 434)| (pix_x == 185 & pix_y == 435)| (pix_x == 185 & pix_y == 436)| (pix_x == 185 & pix_y == 437)| (pix_x == 185 & pix_y == 438)| (pix_x == 186 & pix_y == 206)| (pix_x == 186 & pix_y == 207)| (pix_x == 186 & pix_y == 208)| (pix_x == 186 & pix_y == 251)| (pix_x == 186 & pix_y == 384)| (pix_x == 186 & pix_y == 385)| (pix_x == 186 & pix_y == 432)| (pix_x == 186 & pix_y == 433)| (pix_x == 186 & pix_y == 434)| (pix_x == 186 & pix_y == 435)| (pix_x == 186 & pix_y == 436)| (pix_x == 186 & pix_y == 437)| (pix_x == 186 & pix_y == 438)| (pix_x == 187 & pix_y == 229)| (pix_x == 187 & pix_y == 230)| (pix_x == 187 & pix_y == 271)| (pix_x == 187 & pix_y == 434)| (pix_x == 187 & pix_y == 435)| (pix_x == 187 & pix_y == 436)| (pix_x == 188 & pix_y == 229)| (pix_x == 188 & pix_y == 230)| (pix_x == 188 & pix_y == 271)| (pix_x == 188 & pix_y == 434)| (pix_x == 188 & pix_y == 435)| (pix_x == 188 & pix_y == 436)| (pix_x == 189 & pix_y == 229)| (pix_x == 189 & pix_y == 230)| (pix_x == 189 & pix_y == 271)| (pix_x == 189 & pix_y == 434)| (pix_x == 189 & pix_y == 435)| (pix_x == 189 & pix_y == 436)| (pix_x == 190 & pix_y == 318)| (pix_x == 190 & pix_y == 319)| (pix_x == 190 & pix_y == 355)| (pix_x == 190 & pix_y == 384)| (pix_x == 190 & pix_y == 385)| (pix_x == 191 & pix_y == 318)| (pix_x == 191 & pix_y == 319)| (pix_x == 191 & pix_y == 355)| (pix_x == 191 & pix_y == 384)| (pix_x == 191 & pix_y == 385)| (pix_x == 192 & pix_y == 318)| (pix_x == 192 & pix_y == 319)| (pix_x == 192 & pix_y == 320)| (pix_x == 192 & pix_y == 321)| (pix_x == 192 & pix_y == 427)| (pix_x == 192 & pix_y == 428)| (pix_x == 192 & pix_y == 429)| (pix_x == 192 & pix_y == 430)| (pix_x == 193 & pix_y == 318)| (pix_x == 193 & pix_y == 319)| (pix_x == 193 & pix_y == 320)| (pix_x == 193 & pix_y == 321)| (pix_x == 193 & pix_y == 427)| (pix_x == 193 & pix_y == 428)| (pix_x == 193 & pix_y == 429)| (pix_x == 193 & pix_y == 430)| (pix_x == 194 & pix_y == 407)| (pix_x == 194 & pix_y == 408)| (pix_x == 194 & pix_y == 409)| (pix_x == 194 & pix_y == 410)| (pix_x == 194 & pix_y == 426)| (pix_x == 194 & pix_y == 427)| (pix_x == 194 & pix_y == 428)| (pix_x == 195 & pix_y == 407)| (pix_x == 195 & pix_y == 408)| (pix_x == 195 & pix_y == 409)| (pix_x == 195 & pix_y == 410)| (pix_x == 195 & pix_y == 426)| (pix_x == 195 & pix_y == 427)| (pix_x == 195 & pix_y == 428)| (pix_x == 196 & pix_y == 407)| (pix_x == 196 & pix_y == 408)| (pix_x == 196 & pix_y == 409)| (pix_x == 196 & pix_y == 410)| (pix_x == 196 & pix_y == 426)| (pix_x == 196 & pix_y == 427)| (pix_x == 196 & pix_y == 428)| (pix_x == 197 & pix_y == 373)| (pix_x == 198 & pix_y == 373)| (pix_x == 202 & pix_y == 341)| (pix_x == 202 & pix_y == 342)| (pix_x == 203 & pix_y == 341)| (pix_x == 203 & pix_y == 342)| (pix_x == 204 & pix_y == 340)| (pix_x == 204 & pix_y == 341)| (pix_x == 204 & pix_y == 342)| (pix_x == 204 & pix_y == 381)| (pix_x == 204 & pix_y == 382)| (pix_x == 205 & pix_y == 340)| (pix_x == 205 & pix_y == 341)| (pix_x == 205 & pix_y == 342)| (pix_x == 205 & pix_y == 381)| (pix_x == 205 & pix_y == 382)| (pix_x == 206 & pix_y == 254)| (pix_x == 206 & pix_y == 255)| (pix_x == 206 & pix_y == 259)| (pix_x == 206 & pix_y == 260)| (pix_x == 206 & pix_y == 332)| (pix_x == 206 & pix_y == 340)| (pix_x == 206 & pix_y == 341)| (pix_x == 206 & pix_y == 342)| (pix_x == 206 & pix_y == 355)| (pix_x == 207 & pix_y == 254)| (pix_x == 207 & pix_y == 255)| (pix_x == 207 & pix_y == 259)| (pix_x == 207 & pix_y == 260)| (pix_x == 207 & pix_y == 332)| (pix_x == 207 & pix_y == 340)| (pix_x == 207 & pix_y == 341)| (pix_x == 207 & pix_y == 342)| (pix_x == 207 & pix_y == 355)| (pix_x == 208 & pix_y == 254)| (pix_x == 208 & pix_y == 255)| (pix_x == 208 & pix_y == 259)| (pix_x == 208 & pix_y == 260)| (pix_x == 208 & pix_y == 332)| (pix_x == 208 & pix_y == 340)| (pix_x == 208 & pix_y == 341)| (pix_x == 208 & pix_y == 342)| (pix_x == 208 & pix_y == 355)| (pix_x == 209 & pix_y == 257)| (pix_x == 209 & pix_y == 258)| (pix_x == 209 & pix_y == 259)| (pix_x == 209 & pix_y == 260)| (pix_x == 210 & pix_y == 257)| (pix_x == 210 & pix_y == 258)| (pix_x == 210 & pix_y == 259)| (pix_x == 210 & pix_y == 260)| (pix_x == 214 & pix_y == 242)| (pix_x == 214 & pix_y == 243)| (pix_x == 214 & pix_y == 287)| (pix_x == 214 & pix_y == 288)| (pix_x == 214 & pix_y == 289)| (pix_x == 215 & pix_y == 242)| (pix_x == 215 & pix_y == 243)| (pix_x == 215 & pix_y == 287)| (pix_x == 215 & pix_y == 288)| (pix_x == 215 & pix_y == 289)| (pix_x == 218 & pix_y == 292)| (pix_x == 218 & pix_y == 293)| (pix_x == 219 & pix_y == 292)| (pix_x == 219 & pix_y == 293)| (pix_x == 220 & pix_y == 292)| (pix_x == 220 & pix_y == 293)| (pix_x == 221 & pix_y == 322)| (pix_x == 221 & pix_y == 327)| (pix_x == 221 & pix_y == 356)| (pix_x == 221 & pix_y == 357)| (pix_x == 222 & pix_y == 322)| (pix_x == 222 & pix_y == 327)| (pix_x == 222 & pix_y == 356)| (pix_x == 222 & pix_y == 357)| (pix_x == 223 & pix_y == 322)| (pix_x == 224 & pix_y == 322)| (pix_x == 225 & pix_y == 322)| (pix_x == 226 & pix_y == 264)| (pix_x == 226 & pix_y == 265)| (pix_x == 227 & pix_y == 264)| (pix_x == 227 & pix_y == 265)| (pix_x == 228 & pix_y == 228)| (pix_x == 228 & pix_y == 379)| (pix_x == 228 & pix_y == 380)| (pix_x == 229 & pix_y == 228)| (pix_x == 229 & pix_y == 379)| (pix_x == 229 & pix_y == 380)| (pix_x == 235 & pix_y == 320)| (pix_x == 235 & pix_y == 321)| (pix_x == 235 & pix_y == 330)| (pix_x == 235 & pix_y == 331)| (pix_x == 235 & pix_y == 332)| (pix_x == 236 & pix_y == 320)| (pix_x == 236 & pix_y == 321)| (pix_x == 236 & pix_y == 330)| (pix_x == 236 & pix_y == 331)| (pix_x == 236 & pix_y == 332)| (pix_x == 237 & pix_y == 320)| (pix_x == 237 & pix_y == 321)| (pix_x == 237 & pix_y == 330)| (pix_x == 237 & pix_y == 331)| (pix_x == 237 & pix_y == 332)| (pix_x == 238 & pix_y == 327)| (pix_x == 238 & pix_y == 332)| (pix_x == 239 & pix_y == 327)| (pix_x == 239 & pix_y == 332);
assign win2 = 0;
assign win3 = 0;

//assign win1 = (pix_y > 400) & (pix_y < 450);
//assign win2 = (pix_x > 620) & (pix_x < 630);
//assign win3 = (pix_x > 20) & (pix_x< 640); 
//becomes a 853x480 display on 16:9

assign r_out = win1;
assign g_out = win2;
assign b_out = win3;
//assign temp = win4;

//-----------------------------------------------------------


endmodule
